module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(7), .GND_b_1_row_4(net1920[0:7]), .Vs_b_0_row_4(net124[0:7]), .Vs_b_1_row_4(net125[0:7]), .VINJ_b_1_row_4(net1927[0:7]), .Vsel_b_0_row_4(net1885[0:7]), .Vsel_b_1_row_4(net1886[0:7]), .Vg_b_0_row_4(net1899[0:7]), .Vg_b_1_row_4(net1900[0:7]), .VTUN_brow_4(net1913[0:7]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(17), .matrix_row(5), .matrix_col(9), .GND_b_1_row_4(net285[0:9]), .Vs_b_0_row_4(net286[0:9]), .Vs_b_1_row_4(net287[0:9]), .VINJ_b_1_row_4(net305[0:9]), .Vsel_b_0_row_4(net1964[0:9]), .Vsel_b_1_row_4(net1966[0:9]), .Vg_b_0_row_4(net306[0:9]), .Vg_b_1_row_4(net307[0:9]), .VTUN_brow_4(net308[0:9]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(26), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1940[0:1]), .Vsel_b_0_row_4(net1943[0:1]), .Vsel_b_1_row_4(net1944[0:1]), .Vg_b_0_row_4(net1945[0:1]), .Vg_b_1_row_4(net1946[0:1]), .VTUN_brow_4(net1941[0:1]), .GND_b_1_row_4(net1942[0:1]));
	S_BLOCK_BUFFER I__4 (.island_num(0), .row(0), .col(8), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__5 (.island_num(0), .row(0), .col(9), .matrix_row(4), .matrix_col(1));
	S_BLOCK_CONN_PINS I__6 (.island_num(0), .row(4), .col(9), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__7 (.island_num(0), .row(0), .col(10), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__8 (.island_num(0), .row(3), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__9 (.island_num(0), .row(4), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__10 (.island_num(0), .row(0), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_CONN_PINS I__11 (.island_num(0), .row(2), .col(11), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__12 (.island_num(0), .row(3), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__13 (.island_num(0), .row(0), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_CONN_PINS I__14 (.island_num(0), .row(1), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__15 (.island_num(0), .row(2), .col(12), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__16 (.island_num(0), .row(0), .col(13), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__17 (.island_num(0), .row(1), .col(13), .matrix_row(4), .matrix_col(1));
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1947[0:1]), .Vsel_b_0_row_4(net1950[0:1]), .Vsel_b_1_row_4(net1951[0:1]), .Vg_b_0_row_4(net1952[0:1]), .Vg_b_1_row_4(net1953[0:1]), .VTUN_brow_4(net1948[0:1]), .GND_b_1_row_4(net1949[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1954[0:1]), .Vsel_b_0_row_4(net1957[0:1]), .Vsel_b_1_row_4(net1958[0:1]), .Vg_b_0_row_4(net1959[0:1]), .Vg_b_1_row_4(net1960[0:1]), .VTUN_brow_4(net1955[0:1]), .GND_b_1_row_4(net1956[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(6), .decode_n0_RUN_OUT_0_(net2031), .decode_n0_RUN_OUT_1_(net2032), .decode_n0_RUN_OUT_2_(net2037), .decode_n0_RUN_OUT_3_(net2038), .decode_n1_RUN_OUT_0_(net2043), .decode_n1_RUN_OUT_1_(net2044), .decode_n1_RUN_OUT_2_(net2049), .decode_n1_RUN_OUT_3_(net2050), .decode_n2_RUN_OUT_0_(net2055), .decode_n2_RUN_OUT_1_(net2056), .decode_n2_RUN_OUT_2_(net2061), .decode_n2_RUN_OUT_3_(net2062), .decode_n3_RUN_OUT_0_(net2067), .decode_n3_RUN_OUT_1_(net2068), .decode_n3_RUN_OUT_2_(net2073), .decode_n3_RUN_OUT_3_(net2074), .decode_n4_RUN_OUT_2_(net2079), .decode_n4_RUN_OUT_3_(net2080), .decode_n5_RUN_OUT_0_(net2085), .decode_n5_RUN_OUT_1_(net2086), .decode_n5_RUN_OUT_2_(net2091), .decode_n5_RUN_OUT_3_(net2092), .decode_n6_RUN_OUT_0_(net2097), .decode_n6_RUN_OUT_1_(net2098), .decode_n6_RUN_OUT_2_(net2103), .decode_n6_RUN_OUT_3_(net2104), .decode_n7_RUN_OUT_0_(net2109), .decode_n7_RUN_OUT_1_(net2110), .decode_n7_RUN_OUT_2_(net2115), .decode_n7_RUN_OUT_3_(net2116), .decode_n8_RUN_OUT_0_(net2121), .decode_n8_RUN_OUT_1_(net2122), .decode_n8_RUN_OUT_2_(net2127), .decode_n8_RUN_OUT_3_(net2128), .decode_n9_RUN_OUT_0_(net2133), .decode_n9_RUN_OUT_1_(net2134), .decode_n9_RUN_OUT_2_(net2139), .decode_n9_RUN_OUT_3_(net2140), .decode_n0_OUT_0_(net2029), .decode_n0_OUT_1_(net2030), .decode_n0_OUT_2_(net2035), .decode_n0_OUT_3_(net2036), .decode_n1_OUT_0_(net2041), .decode_n1_OUT_1_(net2042), .decode_n1_OUT_2_(net2047), .decode_n1_OUT_3_(net2048), .decode_n2_OUT_0_(net2053), .decode_n2_OUT_1_(net2054), .decode_n2_OUT_2_(net2059), .decode_n2_OUT_3_(net2060), .decode_n3_OUT_0_(net2065), .decode_n3_OUT_1_(net2066), .decode_n3_OUT_2_(net2071), .decode_n3_OUT_3_(net2072), .decode_n4_OUT_2_(net2077), .decode_n4_OUT_3_(net2078), .decode_n5_OUT_0_(net2083), .decode_n5_OUT_1_(net2084), .decode_n5_OUT_2_(net2089), .decode_n5_OUT_3_(net2090), .decode_n6_OUT_0_(net2095), .decode_n6_OUT_1_(net2096), .decode_n6_OUT_2_(net2101), .decode_n6_OUT_3_(net2102), .decode_n7_OUT_0_(net2107), .decode_n7_OUT_1_(net2108), .decode_n7_OUT_2_(net2113), .decode_n7_OUT_3_(net2114), .decode_n8_OUT_0_(net2119), .decode_n8_OUT_1_(net2120), .decode_n8_OUT_2_(net2125), .decode_n8_OUT_3_(net2126), .decode_n9_OUT_0_(net2131), .decode_n9_OUT_1_(net2132), .decode_n9_OUT_2_(net2137), .decode_n9_OUT_3_(net2138), .decode_n0_VINJ_b_0_(net2027), .decode_n0_VINJ_b_1_(net2033), .decode_n1_VINJ_b_0_(net2039), .decode_n1_VINJ_b_1_(net2045), .decode_n2_VINJ_b_0_(net2051), .decode_n2_VINJ_b_1_(net2057), .decode_n3_VINJ_b_0_(net2063), .decode_n3_VINJ_b_1_(net2069), .decode_n4_VINJ_b_1_(net2075), .decode_n5_VINJ_b_0_(net2081), .decode_n5_VINJ_b_1_(net2087), .decode_n6_VINJ_b_0_(net2093), .decode_n6_VINJ_b_1_(net2099), .decode_n7_VINJ_b_0_(net2105), .decode_n7_VINJ_b_1_(net2111), .decode_n8_VINJ_b_0_(net2117), .decode_n8_VINJ_b_1_(net2123), .decode_n9_VINJ_b_0_(net2129), .decode_n9_VINJ_b_1_(net2135), .decode_n0_GND_b_0_(net2028), .decode_n0_GND_b_1_(net2034), .decode_n1_GND_b_0_(net2040), .decode_n1_GND_b_1_(net2046), .decode_n2_GND_b_0_(net2052), .decode_n2_GND_b_1_(net2058), .decode_n3_GND_b_0_(net2064), .decode_n3_GND_b_1_(net2070), .decode_n4_GND_b_1_(net2076), .decode_n5_GND_b_0_(net2082), .decode_n5_GND_b_1_(net2088), .decode_n6_GND_b_0_(net2094), .decode_n6_GND_b_1_(net2100), .decode_n7_GND_b_0_(net2106), .decode_n7_GND_b_1_(net2112), .decode_n8_GND_b_0_(net2118), .decode_n8_GND_b_1_(net2124), .decode_n9_GND_b_0_(net2130), .decode_n9_GND_b_1_(net2136));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(26), .switch_n0_VPWR_0_(net2031), .switch_n0_VPWR_1_(net2032), .switch_n1_VPWR_0_(net2037), .switch_n1_VPWR_1_(net2038), .switch_n2_VPWR_0_(net2043), .switch_n2_VPWR_1_(net2044), .switch_n3_VPWR_0_(net2049), .switch_n3_VPWR_1_(net2050), .switch_n4_VPWR_0_(net2055), .switch_n4_VPWR_1_(net2056), .switch_n5_VPWR_0_(net2061), .switch_n5_VPWR_1_(net2062), .switch_n6_VPWR_0_(net2067), .switch_n6_VPWR_1_(net2068), .switch_n7_VPWR_0_(net2073), .switch_n7_VPWR_1_(net2074), .switch_n14_VPWR_0_(net2079), .switch_n14_VPWR_1_(net2080), .switch_n16_VPWR_0_(net2085), .switch_n16_VPWR_1_(net2086), .switch_n17_VPWR_0_(net2091), .switch_n17_VPWR_1_(net2092), .switch_n18_VPWR_0_(net2097), .switch_n18_VPWR_1_(net2098), .switch_n19_VPWR_0_(net2103), .switch_n19_VPWR_1_(net2104), .switch_n20_VPWR_0_(net2109), .switch_n20_VPWR_1_(net2110), .switch_n21_VPWR_0_(net2115), .switch_n21_VPWR_1_(net2116), .switch_n22_VPWR_0_(net2121), .switch_n22_VPWR_1_(net2122), .switch_n23_VPWR_0_(net2127), .switch_n23_VPWR_1_(net2128), .switch_n24_VPWR_0_(net2133), .switch_n24_VPWR_1_(net2134), .switch_n25_VPWR_0_(net2139), .switch_n25_VPWR_1_(net2140), .switch_n0_GND_T(net2028), .switch_n1_GND_T(net2034), .switch_n2_GND_T(net2040), .switch_n3_GND_T(net2046), .switch_n4_GND_T(net2052), .switch_n5_GND_T(net2058), .switch_n6_GND_T(net2064), .switch_n7_GND_T(net2070), .switch_n14_GND_T(net2076), .switch_n16_GND_T(net2082), .switch_n17_GND_T(net2088), .switch_n18_GND_T(net2094), .switch_n19_GND_T(net2100), .switch_n20_GND_T(net2106), .switch_n21_GND_T(net2112), .switch_n22_GND_T(net2118), .switch_n23_GND_T(net2124), .switch_n24_GND_T(net2130), .switch_n25_GND_T(net2136), .switch_n0_decode_0_(net2029), .switch_n0_decode_1_(net2030), .switch_n1_decode_0_(net2035), .switch_n1_decode_1_(net2036), .switch_n2_decode_0_(net2041), .switch_n2_decode_1_(net2042), .switch_n3_decode_0_(net2047), .switch_n3_decode_1_(net2048), .switch_n4_decode_0_(net2053), .switch_n4_decode_1_(net2054), .switch_n5_decode_0_(net2059), .switch_n5_decode_1_(net2060), .switch_n6_decode_0_(net2065), .switch_n6_decode_1_(net2066), .switch_n7_decode_0_(net2071), .switch_n7_decode_1_(net2072), .switch_n14_decode_0_(net2077), .switch_n14_decode_1_(net2078), .switch_n16_decode_0_(net2083), .switch_n16_decode_1_(net2084), .switch_n17_decode_0_(net2089), .switch_n17_decode_1_(net2090), .switch_n18_decode_0_(net2095), .switch_n18_decode_1_(net2096), .switch_n19_decode_0_(net2101), .switch_n19_decode_1_(net2102), .switch_n20_decode_0_(net2107), .switch_n20_decode_1_(net2108), .switch_n21_decode_0_(net2113), .switch_n21_decode_1_(net2114), .switch_n22_decode_0_(net2119), .switch_n22_decode_1_(net2120), .switch_n23_decode_0_(net2125), .switch_n23_decode_1_(net2126), .switch_n24_decode_0_(net2131), .switch_n24_decode_1_(net2132), .switch_n25_decode_0_(net2137), .switch_n25_decode_1_(net2138), .switch_n0_VINJ_T(net2027), .switch_n1_VINJ_T(net2033), .switch_n2_VINJ_T(net2039), .switch_n3_VINJ_T(net2045), .switch_n4_VINJ_T(net2051), .switch_n5_VINJ_T(net2057), .switch_n6_VINJ_T(net2063), .switch_n7_VINJ_T(net2069), .switch_n14_VINJ_T(net2075), .switch_n16_VINJ_T(net2081), .switch_n17_VINJ_T(net2087), .switch_n18_VINJ_T(net2093), .switch_n19_VINJ_T(net2099), .switch_n20_VINJ_T(net2105), .switch_n21_VINJ_T(net2111), .switch_n22_VINJ_T(net2117), .switch_n23_VINJ_T(net2123), .switch_n24_VINJ_T(net2129), .switch_n25_VINJ_T(net2135));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch));
	none switch_ind(.island_num(0), .direction(horizontal), .col(8));
	none switch_ind(.island_num(0), .direction(horizontal), .col(9));
	none switch_ind(.island_num(0), .direction(horizontal), .col(10));
	none switch_ind(.island_num(0), .direction(horizontal), .col(11));
	none switch_ind(.island_num(0), .direction(horizontal), .col(12));
	none switch_ind(.island_num(0), .direction(horizontal), .col(13));
	none switch_ind(.island_num(0), .direction(horizontal), .col(15));


	/* Island 1 */
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__0 (.island_num(1), .row(0), .col(0), .matrix_row(1), .matrix_col(8));
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(7), .matrix_col(8), .GND_b_0_row_6(net1109[0:8]), .GND_b_1_row_6(net1110[0:8]), .Vs_b_0_row_6(net1119[0:8]), .Vs_b_1_row_6(net1120[0:8]), .VINJ_b_0_row_6(net1123[0:8]), .VINJ_b_1_row_6(net1124[0:8]), .Vsel_b_0_row_6(net1127[0:8]), .Vsel_b_1_row_6(net1128[0:8]), .Vg_b_0_row_6(net1131[0:8]), .Vg_b_1_row_6(net1132[0:8]), .VTUN_brow_6(net1135[0:8]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(8), .matrix_row(6), .matrix_col(10));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(7), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1784), .P_1_row_0(net1785), .A_0_row_0(net1786), .A_1_row_0(net1787), .A_2_row_0(net1788), .A_3_row_0(net1789));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1797), .P_1_row_0(net1798), .A_0_row_0(net1799), .A_1_row_0(net1800), .A_2_row_0(net1801), .A_3_row_0(net1802));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1815), .P_1_row_0(net1816), .A_0_row_0(net1817), .A_1_row_0(net1818), .A_2_row_0(net1819), .A_3_row_0(net1820));
	TSMC350nm_4TGate_ST_BMatrix_NoSwitch I__8 (.island_num(1), .row(3), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1833), .P_1_row_0(net1834), .P_2_row_0(net1835), .P_3_row_0(net1836), .A_0_row_0(net1837), .A_1_row_0(net1838), .A_2_row_0(net1839), .A_3_row_0(net1840));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1852), .P_1_row_0(net1853), .P_2_row_0(net1854), .P_3_row_0(net1855), .A_0_row_0(net1856), .A_1_row_0(net1857));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1867), .A_1_row_0(net1868), .A_2_row_0(net1869), .A_3_row_0(net1870));
	TSMC350nm_4TGate_ST_BMatrix I__11 (.island_num(1), .row(6), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1875), .A_1_row_0(net1876), .A_2_row_0(net1877), .A_3_row_0(net1878));
	TSMC350nm_4TGate_ST_BMatrix I__12 (.island_num(1), .row(7), .col(18), .matrix_row(1), .matrix_col(1));
	TSMC350nm_OutMtrx_IndrctSwcs I__13 (.island_num(1), .row(9), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__14 (.island_num(1), .row(10), .col(8), .matrix_row(2), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__15 (.island_num(1), .row(10), .col(18), .matrix_row(2), .matrix_col(1));
	TSMC350nm_TA2Cell_Weak cab_device_16 (.island_num(1), .row(2), .col(19), .VD_P_0_(net1784), .VD_P_1_(net1785), .VIN1_PLUS(net1786), .VIN1_MINUS(net1787), .VIN2_PLUS(net1788), .VIN2_MINUS(net1789), .OUTPUT_0_(net1790[0]), .OUTPUT_1_(net1791[0]), .Vsel_0_(net1861), .Vsel_1_(net1862), .RUN(net1792), .Vg_0_(net1863), .Vg_1_(net1864), .PROG(net1793), .VTUN(net1794), .VINJ(net1795), .GND(net1796), .VPWR(net1873), .Vsel_b_0_(net1805), .Vsel_b_1_(net1806), .RUN_b(net1807), .Vg_b_0_(net1808), .Vg_b_1_(net1809), .PROG_b(net1810), .VTUN_b(net1811), .VINJ_b(net1812), .GND_b(net1813), .VPWR_b(net1814));
	TSMC350nm_TA2Cell_Weak cab_device_17 (.island_num(1), .row(3), .col(19), .VD_P_0_(net1797), .VD_P_1_(net1798), .VIN1_PLUS(net1799), .VIN1_MINUS(net1800), .VIN2_PLUS(net1801), .VIN2_MINUS(net1802), .OUTPUT_0_(net1803[0]), .OUTPUT_1_(net1804[0]), .Vsel_0_(net1805), .Vsel_1_(net1806), .RUN(net1807), .Vg_0_(net1808), .Vg_1_(net1809), .PROG(net1810), .VTUN(net1811), .VINJ(net1812), .GND(net1813), .VPWR(net1814), .Vsel_b_0_(net1823), .Vsel_b_1_(net1824), .RUN_b(net1825), .Vg_b_0_(net1826), .Vg_b_1_(net1827), .PROG_b(net1828), .VTUN_b(net1829), .VINJ_b(net1830), .GND_b(net1831), .VPWR_b(net1832));
	TSMC350nm_TA2Cell_Strong cab_device_18 (.island_num(1), .row(4), .col(19), .VD_P_0_(net1815), .VD_P_1_(net1816), .VIN1_PLUS(net1817), .VIN1_MINUS(net1818), .VIN2_PLUS(net1819), .VIN2_MINUS(net1820), .OUTPUT_0_(net1821[0]), .OUTPUT_1_(net1822[0]), .Vsel_0_(net1823), .Vsel_1_(net1824), .RUN(net1825), .Vg_0_(net1826), .Vg_1_(net1827), .PROG(net1828), .VTUN(net1829), .VINJ(net1830), .GND(net1831), .VPWR(net1832), .Vg_b_0_(net1848), .PROG_b(net1851), .VTUN_b(net1849), .VINJ_b(net1847), .GND_b(net1850));
	TSMC350nm_4WTA_IndirectProg cab_device_19 (.island_num(1), .row(5), .col(19), .VD_P_0_(net1833), .VD_P_1_(net1834), .VD_P_2_(net1835), .VD_P_3_(net1836), .Iin_0_(net1837), .Iin_1_(net1838), .Iin_2_(net1839), .Iin_3_(net1840), .Vout_0_(net1841[0]), .Vout_1_(net1842[0]), .Vout_2_(net1843[0]), .Vout_3_(net1844[0]), .Vmid(net1845[0]), .Vbias(net1846[0]), .Vsel(net1861), .Vs(net1873), .VINJ(net1847), .Vg(net1848), .VTUN(net1849), .GND(net1850), .PROG(net1851), .VINJ_b(net1860), .VTUN_b(net1866), .GND_b(net1865));
	TSMC350nm_Cap_Bank cab_device_20 (.island_num(1), .row(6), .col(19), .VD_P_0_(net1852), .VD_P_1_(net1853), .VD_P_2_(net1854), .VD_P_3_(net1855), .VIN_0_(net1856), .VIN_1_(net1857), .OUT_0_(net1858[0]), .OUT_1_(net1859[0]), .VINJ(net1860), .Vsel_0_(net1861), .Vsel_1_(net1862), .Vg_0_(net1863), .Vg_1_(net1864), .GND(net1865), .VTUN(net1866), .GND_b(net1874));
	TSMC350nm_NandPfets cab_device_21 (.island_num(1), .row(7), .col(19), .GATE_N(net1867), .SOURCE_N(net1868), .GATE_P(net1869), .SOURCE_P(net1870), .DRAIN_N(net1871[0]), .DRAIN_P(net1872[0]), .VPWR(net1873), .GND(net1874), .VPWR_b(net1882), .GND_b(net1883));
	TSMC350nm_TGate_2nMirror cab_device_22 (.island_num(1), .row(8), .col(19), .IN_CM_0_(net1875), .IN_CM_1_(net1876), .SelN(net1877), .IN_TG(net1878), .OUT_CM_0_(net1879[0]), .OUT_CM_1_(net1880[0]), .OUT_TG(net1881[0]), .VPWR(net1882), .GND(net1883));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(1), .direction(vertical), .num(12), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(12), .type(prog_switch));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(20), .switch_n0_Input_0_(net1884), .switch_n0_Input_1_(net1920[0]), .switch_n1_Input_0_(net124[1]), .switch_n1_Input_1_(net125[1]), .switch_n2_Input_0_(net124[2]), .switch_n2_Input_1_(net125[2]), .switch_n3_Input_0_(net124[3]), .switch_n3_Input_1_(net125[3]), .switch_n4_Input_0_(net286[0]), .switch_n4_Input_1_(net287[0]), .switch_n5_Input_0_(net286[1]), .switch_n5_Input_1_(net287[1]), .switch_n6_Input_0_(net286[2]), .switch_n6_Input_1_(net287[2]), .switch_n7_Input_0_(net286[3]), .switch_n7_Input_1_(net287[3]), .switch_n8_Input_0_(net2203[0]), .switch_n8_Input_1_(net1790[0]), .switch_n9_Input_0_(net1791[0]), .switch_n9_Input_1_(net1803[0]), .switch_n10_Input_0_(net1804[0]), .switch_n10_Input_1_(net1821[0]), .switch_n11_Input_0_(net1822[0]), .switch_n11_Input_1_(net1841[0]), .switch_n12_Input_0_(net1842[0]), .switch_n12_Input_1_(net1843[0]), .switch_n13_Input_0_(net1844[0]), .switch_n13_Input_1_(net1845[0]), .switch_n14_Input_0_(net1846[0]), .switch_n14_Input_1_(net1858[0]), .switch_n15_Input_0_(net1859[0]), .switch_n15_Input_1_(net1871[0]), .switch_n16_Input_0_(net1872[0]), .switch_n16_Input_1_(net1879[0]), .switch_n17_Input_0_(net1880[0]), .switch_n17_Input_1_(net1881[0]), .switch_n0_GND(net1920[0]), .switch_n1_GND(net1920[1]), .switch_n2_GND(net1920[2]), .switch_n3_GND(net1920[3]), .switch_n4_GND(net1920[4]), .switch_n5_GND(net1920[5]), .switch_n6_GND(net1920[6]), .switch_n7_GND(net1942[0]), .switch_n8_GND(net1949[0]), .switch_n9_GND(net1956[0]), .switch_n10_GND(net285[0]), .switch_n11_GND(net285[1]), .switch_n12_GND(net285[2]), .switch_n13_GND(net285[3]), .switch_n14_GND(net285[4]), .switch_n15_GND(net285[5]), .switch_n16_GND(net285[6]), .switch_n17_GND(net285[7]), .switch_n0_Vsel_0_(net1885[0]), .switch_n0_Vsel_1_(net1886[0]), .switch_n1_Vsel_0_(net1885[1]), .switch_n1_Vsel_1_(net1886[1]), .switch_n2_Vsel_0_(net1885[2]), .switch_n2_Vsel_1_(net1886[2]), .switch_n3_Vsel_0_(net1885[3]), .switch_n3_Vsel_1_(net1886[3]), .switch_n4_Vsel_0_(net1885[4]), .switch_n4_Vsel_1_(net1886[4]), .switch_n5_Vsel_0_(net1885[5]), .switch_n5_Vsel_1_(net1886[5]), .switch_n6_Vsel_0_(net1885[6]), .switch_n6_Vsel_1_(net1886[6]), .switch_n7_Vsel_0_(net1944[0]), .switch_n7_Vsel_1_(net1943[0]), .switch_n8_Vsel_0_(net1951[0]), .switch_n8_Vsel_1_(net1950[0]), .switch_n9_Vsel_0_(net1958[0]), .switch_n9_Vsel_1_(net1957[0]), .switch_n10_Vsel_0_(net1964[0]), .switch_n10_Vsel_1_(net1966[0]), .switch_n11_Vsel_0_(net1964[1]), .switch_n11_Vsel_1_(net1966[1]), .switch_n12_Vsel_0_(net1964[2]), .switch_n12_Vsel_1_(net1966[2]), .switch_n13_Vsel_0_(net1964[3]), .switch_n13_Vsel_1_(net1966[3]), .switch_n14_Vsel_0_(net1964[4]), .switch_n14_Vsel_1_(net1966[4]), .switch_n15_Vsel_0_(net1964[5]), .switch_n15_Vsel_1_(net1966[5]), .switch_n16_Vsel_0_(net1964[6]), .switch_n16_Vsel_1_(net1966[6]), .switch_n17_Vsel_0_(net1964[7]), .switch_n17_Vsel_1_(net1966[7]), .switch_n0_Vg_global_0_(net1899[0]), .switch_n0_Vg_global_1_(net1900[0]), .switch_n1_Vg_global_0_(net1899[1]), .switch_n1_Vg_global_1_(net1900[1]), .switch_n2_Vg_global_0_(net1899[2]), .switch_n2_Vg_global_1_(net1900[2]), .switch_n3_Vg_global_0_(net1899[3]), .switch_n3_Vg_global_1_(net1900[3]), .switch_n4_Vg_global_0_(net1899[4]), .switch_n4_Vg_global_1_(net1900[4]), .switch_n5_Vg_global_0_(net1899[5]), .switch_n5_Vg_global_1_(net1900[5]), .switch_n6_Vg_global_0_(net1899[6]), .switch_n6_Vg_global_1_(net1900[6]), .switch_n7_Vg_global_0_(net1946[0]), .switch_n7_Vg_global_1_(net1945[0]), .switch_n8_Vg_global_0_(net1953[0]), .switch_n8_Vg_global_1_(net1952[0]), .switch_n9_Vg_global_0_(net1960[0]), .switch_n9_Vg_global_1_(net1959[0]), .switch_n10_Vg_global_0_(net306[0]), .switch_n10_Vg_global_1_(net307[0]), .switch_n11_Vg_global_0_(net306[1]), .switch_n11_Vg_global_1_(net307[1]), .switch_n12_Vg_global_0_(net306[2]), .switch_n12_Vg_global_1_(net307[2]), .switch_n13_Vg_global_0_(net306[3]), .switch_n13_Vg_global_1_(net307[3]), .switch_n14_Vg_global_0_(net306[4]), .switch_n14_Vg_global_1_(net307[4]), .switch_n15_Vg_global_0_(net306[5]), .switch_n15_Vg_global_1_(net307[5]), .switch_n16_Vg_global_0_(net306[6]), .switch_n16_Vg_global_1_(net307[6]), .switch_n17_Vg_global_0_(net306[7]), .switch_n17_Vg_global_1_(net307[7]), .switch_n0_VTUN(net1913[0]), .switch_n1_VTUN(net1913[1]), .switch_n2_VTUN(net1913[2]), .switch_n3_VTUN(net1913[3]), .switch_n4_VTUN(net1913[4]), .switch_n5_VTUN(net1913[5]), .switch_n6_VTUN(net1913[6]), .switch_n7_VTUN(net1941[0]), .switch_n8_VTUN(net1948[0]), .switch_n9_VTUN(net1955[0]), .switch_n10_VTUN(net308[0]), .switch_n11_VTUN(net308[1]), .switch_n12_VTUN(net308[2]), .switch_n13_VTUN(net308[3]), .switch_n14_VTUN(net308[4]), .switch_n15_VTUN(net308[5]), .switch_n16_VTUN(net308[6]), .switch_n17_VTUN(net308[7]), .switch_n0_VINJ(net1927[0]), .switch_n1_VINJ(net1927[1]), .switch_n2_VINJ(net1927[2]), .switch_n3_VINJ(net1927[3]), .switch_n4_VINJ(net1927[4]), .switch_n5_VINJ(net1927[5]), .switch_n6_VINJ(net1927[6]), .switch_n7_VINJ(net1940[0]), .switch_n8_VINJ(net1947[0]), .switch_n9_VINJ(net1954[0]), .switch_n10_VINJ(net305[0]), .switch_n11_VINJ(net305[1]), .switch_n12_VINJ(net305[2]), .switch_n13_VINJ(net305[3]), .switch_n14_VINJ(net305[4]), .switch_n15_VINJ(net305[5]), .switch_n16_VINJ(net305[6]), .switch_n17_VINJ(net305[7]));
	none switch_ind(.island_num(1), .direction(horizontal), .col(18));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(19), .VPWR_0_(net1884), .VPWR_1_(net1884), .decode_0_(net1964[8]), .decode_1_(net1966[8]), .GND(net1796), .CTRL_B_0_(net1861), .CTRL_B_1_(net1862), .run_r(net1792), .prog_r(net1793), .Vg_0_(net1863), .Vg_1_(net1864), .VTUN(net1794), .VINJ(net1795), .VDD_1_(net1873));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net1119[0:6]), .out_1_row_0(net1120[0:6]), .VINJ_0_row_0(net1123[0:6]), .VINJ_1_row_0(net1124[0:6]), .Vsel_0_row_0(net1127[0:6]), .Vsel_1_row_0(net1128[0:6]), .Vg_0_row_0(net1131[0:6]), .Vg_1_row_0(net1132[0:6]), .GNDrow_0(net1109[0:6]), .VTUNrow_0(net1135[0:6]), .Dcol_0(net124[6:7]), .CLKcol_0(net125[6:7]), .Qcol_5(net125[6:7]), .comcol_0(net2203[0:1]));

 	/*Programming Mux */ 

 endmodule