VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  CAPACITANCE PICOFARADS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER OD
  TYPE MASTERSLICE ;
END OD

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER PP
  TYPE IMPLANT ;
  WIDTH 0.18 ;
  SPACING 0.18 ;
  AREA 0.122 ;
END PP

LAYER NP
  TYPE IMPLANT ;
  WIDTH 0.18 ;
  SPACING 0.18 ;
  AREA 0.122 ;
END NP

LAYER CO
  TYPE CUT ;
  SPACING 0.11 ;
  SPACING 0.11 ;
  SPACING 0.12 ;
  SPACING 0.14 ADJACENTCUTS 3 WITHIN 0.15 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 10 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 10 ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.18 ;
  WIDTH 0.09 ;
  OFFSET 0.09 ;
  AREA 0.042 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 0.384 0.424 1.504 4.504 
    WIDTH 0.004 0.09 0.09 0.09 0.09 0.09 
    WIDTH 0.204 0.09 0.11 0.09 0.09 0.09 
    WIDTH 0.424 0.09 0.11 0.16 0.09 0.09 
    WIDTH 1.504 0.09 0.11 0.16 0.5 0.09 
    WIDTH 4.504 0.09 0.11 0.16 0.5 1.5 ;
  MINIMUMCUT 1 WIDTH 0.089 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.099 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.299 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 0.699 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.0868 ;
  CAPACITANCE CPERSQDIST 0.00514 ;
  THICKNESS 1800 ;
  EDGECAPACITANCE 0.00758 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       9.36775 19.5501 39.9148 80.6441 253.744 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       1.20706 2.15515 3.93091 7.39472 21.9815 ;
END M1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 0.384 0.404 1.504 4.504 
    WIDTH 0.004 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.204 0.1 0.12 0.1 0.1 0.1 
    WIDTH 0.404 0.1 0.12 0.16 0.1 0.1 
    WIDTH 1.504 0.1 0.12 0.16 0.5 0.1 
    WIDTH 4.504 0.1 0.12 0.16 0.5 1.5 ;
  MINIMUMCUT 1 WIDTH 0.089 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.099 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 4 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.00298 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00659 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.749923 1.31913 2.37142 4.41089 12.9754 ;
END M2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 0.384 0.404 1.504 4.504 
    WIDTH 0.004 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.204 0.1 0.12 0.1 0.1 0.1 
    WIDTH 0.404 0.1 0.12 0.16 0.1 0.1 
    WIDTH 1.504 0.1 0.12 0.16 0.5 0.1 
    WIDTH 4.504 0.1 0.12 0.16 0.5 1.5 ;
  MINIMUMCUT 1 WIDTH 0.099 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 4 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.00199 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00578 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.696634 1.16947 1.99669 3.54867 9.95791 ;
END M3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 0.384 0.404 1.504 4.504 
    WIDTH 0.004 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.204 0.1 0.12 0.1 0.1 0.1 
    WIDTH 0.404 0.1 0.12 0.16 0.1 0.1 
    WIDTH 1.504 0.1 0.12 0.16 0.5 0.1 
    WIDTH 4.504 0.1 0.12 0.16 0.5 1.5 ;
  MINIMUMCUT 1 WIDTH 0.099 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 4 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.00149 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00537 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.674844 1.10631 1.83204 3.15479 8.51792 ;
END M4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 0.384 0.404 1.504 4.504 
    WIDTH 0.004 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.204 0.1 0.12 0.1 0.1 0.1 
    WIDTH 0.404 0.1 0.12 0.16 0.1 0.1 
    WIDTH 1.504 0.1 0.12 0.16 0.5 0.1 
    WIDTH 4.504 0.1 0.12 0.16 0.5 1.5 ;
  MINIMUMCUT 1 WIDTH 0.099 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 4 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.0012 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00513 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.59004 0.967284 1.60182 2.75834 7.44752 ;
END M5

LAYER VIA5
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 0.384 0.404 1.504 4.504 
    WIDTH 0.004 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.204 0.1 0.12 0.1 0.1 0.1 
    WIDTH 0.404 0.1 0.12 0.16 0.1 0.1 
    WIDTH 1.504 0.1 0.12 0.16 0.5 0.1 
    WIDTH 4.504 0.1 0.12 0.16 0.5 1.5 ;
  MINIMUMCUT 1 WIDTH 0.099 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 4 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.000996 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00502 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.531302 0.870991 1.44236 2.48375 6.70612 ;
END M6

LAYER VIA6
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 0.384 0.404 1.504 4.504 
    WIDTH 0.004 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.204 0.1 0.12 0.1 0.1 0.1 
    WIDTH 0.404 0.1 0.12 0.16 0.1 0.1 
    WIDTH 1.504 0.1 0.12 0.16 0.5 0.1 
    WIDTH 4.504 0.1 0.12 0.16 0.5 1.5 ;
  MINIMUMCUT 1 WIDTH 0.099 ;
  MINIMUMCUT 2 WIDTH 0.299 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.699 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.359 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.799 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 1.8 FROMABOVE LENGTH 1.8 WITHIN 1.7 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.000854 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00529 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.486946 0.798276 1.32194 2.2764 6.14627 ;
END M7

LAYER VIA7
  TYPE CUT ;
  SPACING 0.34 ;
  SPACING 0.34 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.8 ;
  WIDTH 0.4 ;
  OFFSET 0.4 ;
  AREA 0.565 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 1.504 4.504 
    WIDTH 0.004 0.4 0.4 0.4 
    WIDTH 1.504 0.4 0.5 0.5 
    WIDTH 4.504 0.4 0.5 1.5 ;
  MINIMUMCUT 1 WIDTH 0.099 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.359 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.799 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.359 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.8 FROMBELOW LENGTH 1.8 WITHIN 1.7 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 1.8 FROMABOVE LENGTH 1.8 WITHIN 1.7 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.565 ;
  RESISTANCE RPERSQ 0.0215 ;
  CAPACITANCE CPERSQDIST 0.00323 ;
  THICKNESS 9000 ;
  EDGECAPACITANCE 0.00615 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       16.0372 33.8563 69.4945 140.771 443.695 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       1.29043 2.05444 3.2317 5.20772 12.6666 ;
END M8

LAYER VIA8
  TYPE CUT ;
  SPACING 0.34 ;
  SPACING 0.34 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 4 ;
  WIDTH 2 ;
  OFFSET 2 ;
  AREA 9 ;
  SPACING 2 ;
  MINIMUMCUT 2 WIDTH 0.359 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.8 FROMBELOW LENGTH 1.8 WITHIN 1.7 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 9 ;
  RESISTANCE RPERSQ 0.0215 ;
  CAPACITANCE CPERSQDIST 0.00245 ;
  THICKNESS 34000 ;
  EDGECAPACITANCE 0.00564 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 80 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       16.0372 33.8563 69.4945 140.771 443.695 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       1.64281 2.60223 4.05931 6.46339 15.3636 ;
END M9

LAYER RV
  TYPE CUT ;
  SPACING 3 ;
END RV

LAYER AP
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 3 ;
  SPACING 2 ;
  MAXWIDTH 35 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 70 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
END AP

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

MAXVIASTACK 4 RANGE M1 M7 ;
VIARULE AP_M9 GENERATE
  LAYER M9 ;
    ENCLOSURE 1.5 1.5 ;
  LAYER AP ;
    ENCLOSURE 1.5 1.5 ;
  LAYER RV ;
    RECT -1.5 -1.5 1.5 1.5 ;
    SPACING 6 BY 6 ;
END AP_M9

VIARULE M9_M8 GENERATE
  LAYER M8 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER M9 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.7 BY 0.7 ;
END M9_M8

VIARULE M8_M7 GENERATE
  LAYER M7 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER M8 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER VIA7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.7 BY 0.7 ;
END M8_M7

VIARULE M7_M6 GENERATE
  LAYER M6 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M7 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M7_M6

VIARULE M6_M5 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M6 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M6_M5

VIARULE M5_M4 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M5 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M5_M4

VIARULE M4_M3 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M4 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M2_M1

VIARULE M1_PO GENERATE
  LAYER PO ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_PO

VIARULE M1_NPO GENERATE
  LAYER PO ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_NPO

VIARULE M1_PPO GENERATE
  LAYER PO ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_PPO

VIARULE M1_OD GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_OD

VIARULE M1_NOD GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_NOD

VIARULE M1_POD GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_POD

VIARULE M1_NW GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_NW

VIARULE M1_SUB GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_SUB

VIA DFM_M7_M6s
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M6 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M7_M6s

VIA DFM_M6_M5s
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M5 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M6_M5s

VIA DFM_M5_M4s
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M4 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M5_M4s

VIA DFM_M4_M3s
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M3 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M4_M3s

VIA DFM_M3_M2s
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M2 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M3_M2s

VIA DFM_M2_M1s
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M1 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M2_M1s

VIA DFM_M1_ODs
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M1 ;
    RECT -0.105 -0.105 0.105 0.105 ;
  LAYER OD ;
    RECT -0.085 -0.085 0.085 0.085 ;
END DFM_M1_ODs

VIA DFM_M1_POs
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M1 ;
    RECT -0.105 -0.105 0.105 0.105 ;
  LAYER PO ;
    RECT -0.105 -0.105 0.105 0.105 ;
END DFM_M1_POs

VIA AP_M9s
  LAYER RV ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER AP ;
    RECT -3 -3 3 3 ;
  LAYER M9 ;
    RECT -3 -3 3 3 ;
END AP_M9s

VIA M9_M8s
  LAYER VIA8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M9 ;
    RECT -0.58 -0.58 0.58 0.58 ;
  LAYER M8 ;
    RECT -0.26 -0.26 0.26 0.26 ;
END M9_M8s

VIA M8_M7s
  LAYER VIA7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M8 ;
    RECT -0.26 -0.26 0.26 0.26 ;
  LAYER M7 ;
    RECT -0.26 -0.26 0.26 0.26 ;
END M8_M7s

VIA M7_M6s
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M6 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M7_M6s

VIA M6_M5s
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M5 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M6_M5s

VIA M5_M4s
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M4 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M5_M4s

VIA M4_M3s
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M3 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M4_M3s

VIA M3_M2s
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M2 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M3_M2s

VIA M2_M1s
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M1 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M2_M1s

VIA M1_ODs
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER OD ;
    RECT -0.075 -0.075 0.075 0.075 ;
END M1_ODs

VIA M1_POs
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER PO ;
    RECT -0.085 -0.085 0.085 0.085 ;
END M1_POs

VIA M2_M1c
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M1 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M2 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M2_M1c

VIA M3_M2c
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M3 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M3_M2c

VIA M4_M3c
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M4 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M4_M3c

VIA M5_M4c
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M5 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M5_M4c

VIA M6_M5c
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M6 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M6_M5c

VIA M7_M6c
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M7 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M7_M6c

VIA M8_M7c
  LAYER VIA7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M7 ;
    RECT -0.2 -0.26 0.2 0.26 ;
  LAYER M8 ;
    RECT -0.26 -0.2 0.26 0.2 ;
END M8_M7c

VIA M9_M8c
  LAYER VIA8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M8 ;
    RECT -0.48 -0.26 0.48 0.26 ;
  LAYER M9 ;
    RECT -0.26 -0.48 0.26 0.48 ;
END M9_M8c

VIA AP_M9c
  LAYER RV ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER M9 ;
    RECT -3 -3 3 3 ;
  LAYER AP ;
    RECT -3 -3 3 3 ;
END AP_M9c

VIA DFM_M2_M1c
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M1 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M2 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M2_M1c

VIA DFM_M3_M2c
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M3 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M3_M2c

VIA DFM_M4_M3c
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M4 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M4_M3c

VIA DFM_M5_M4c
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M5 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M5_M4c

VIA DFM_M6_M5c
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M6 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M6_M5c

VIA DFM_M7_M6c
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M7 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M7_M6c

SPACING
  SAMENET PO PO 0.12 ;
  SAMENET M1 M1 0.09 ;
  SAMENET M2 M2 0.1 ;
  SAMENET M3 M3 0.1 ;
  SAMENET M4 M4 0.1 ;
  SAMENET M5 M5 0.1 ;
  SAMENET M6 M6 0.1 ;
  SAMENET M7 M7 0.1 ;
  SAMENET M8 M8 0.4 ;
  SAMENET M9 M9 2 ;
  SAMENET VIA1 CO 0 ;
  SAMENET VIA2 VIA1 0 STACK ;
  SAMENET VIA3 VIA2 0 STACK ;
  SAMENET VIA4 VIA3 0 STACK ;
  SAMENET VIA5 VIA4 0 STACK ;
  SAMENET VIA6 VIA5 0 STACK ;
  SAMENET VIA7 VIA6 0 STACK ;
  SAMENET VIA8 VIA7 0 ;
END SPACING

NONDEFAULTRULE LEFDefaultRouteSpec_DFM
  LAYER M9
    WIDTH 2 ;
  END M9
  LAYER M8
    WIDTH 0.4 ;
  END M8
  LAYER M7
    WIDTH 0.1 ;
  END M7
  LAYER M6
    WIDTH 0.1 ;
  END M6
  LAYER M5
    WIDTH 0.1 ;
  END M5
  LAYER M4
    WIDTH 0.1 ;
  END M4
  LAYER M3
    WIDTH 0.1 ;
  END M3
  LAYER M2
    WIDTH 0.1 ;
  END M2
  LAYER M1
    WIDTH 0.09 ;
  END M1
  LAYER PO
    WIDTH 0.06 ;
  END PO
END LEFDefaultRouteSpec_DFM