module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(16), .matrix_col(32), .Vd_R_0_col_32(net1482[0:16]),.Vd_R_1_col_32(net1483[0:16]),.Vd_R_2_col_32(net1484[0:16]),.Vd_R_3_col_32(net1485[0:16]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(6));
	TSMC350nm_GateMuxSwcTile switch(.island_num(0), .direction(horizontal), .num(32));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect01d3 switch(.island_num(0), .direction(vertical), .num(16), .type(drain_select));
	TSMC350nm_FourTgate_ThickOx_FG_MEM switch(.island_num(0), .direction(vertical), .num(16), .type(prog_switch));


	/* Island 1 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(1), .row(0), .col(0), .matrix_row(16), .matrix_col(32));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(1), .direction(horizontal), .bits(6), .decode_n0_VGRUN_0_(net1482[0]),.decode_n0_VGRUN_1_(net1483[0]),.decode_n0_VGRUN_2_(net1484[0]),.decode_n0_VGRUN_3_(net1485[0]),.decode_n1_VGRUN_0_(net1482[1]),.decode_n1_VGRUN_1_(net1483[1]),.decode_n1_VGRUN_2_(net1484[1]),.decode_n1_VGRUN_3_(net1485[1]),.decode_n2_VGRUN_0_(net1482[2]),.decode_n2_VGRUN_1_(net1483[2]),.decode_n2_VGRUN_2_(net1484[2]),.decode_n2_VGRUN_3_(net1485[2]),.decode_n3_VGRUN_0_(net1482[3]),.decode_n3_VGRUN_1_(net1483[3]),.decode_n3_VGRUN_2_(net1484[3]),.decode_n3_VGRUN_3_(net1485[3]),.decode_n4_VGRUN_0_(net1482[4]),.decode_n4_VGRUN_1_(net1483[4]),.decode_n4_VGRUN_2_(net1484[4]),.decode_n4_VGRUN_3_(net1485[4]),.decode_n5_VGRUN_0_(net1482[5]),.decode_n5_VGRUN_1_(net1483[5]),.decode_n5_VGRUN_2_(net1484[5]),.decode_n5_VGRUN_3_(net1485[5]),.decode_n6_VGRUN_0_(net1482[6]),.decode_n6_VGRUN_1_(net1483[6]),.decode_n6_VGRUN_2_(net1484[6]),.decode_n6_VGRUN_3_(net1485[6]),.decode_n7_VGRUN_0_(net1482[7]),.decode_n7_VGRUN_1_(net1483[7]),.decode_n7_VGRUN_2_(net1484[7]),.decode_n7_VGRUN_3_(net1485[7]),.decode_n8_VGRUN_0_(net1482[8]),.decode_n8_VGRUN_1_(net1483[8]),.decode_n8_VGRUN_2_(net1484[8]),.decode_n8_VGRUN_3_(net1485[8]),.decode_n9_VGRUN_0_(net1482[9]),.decode_n9_VGRUN_1_(net1483[9]),.decode_n9_VGRUN_2_(net1484[9]),.decode_n9_VGRUN_3_(net1485[9]),.decode_n10_VGRUN_0_(net1482[10]),.decode_n10_VGRUN_1_(net1483[10]),.decode_n10_VGRUN_2_(net1484[10]),.decode_n10_VGRUN_3_(net1485[10]),.decode_n11_VGRUN_0_(net1482[11]),.decode_n11_VGRUN_1_(net1483[11]),.decode_n11_VGRUN_2_(net1484[11]),.decode_n11_VGRUN_3_(net1485[11]),.decode_n12_VGRUN_0_(net1482[12]),.decode_n12_VGRUN_1_(net1483[12]),.decode_n12_VGRUN_2_(net1484[12]),.decode_n12_VGRUN_3_(net1485[12]),.decode_n13_VGRUN_0_(net1482[13]),.decode_n13_VGRUN_1_(net1483[13]),.decode_n13_VGRUN_2_(net1484[13]),.decode_n13_VGRUN_3_(net1485[13]),.decode_n14_VGRUN_0_(net1482[14]),.decode_n14_VGRUN_1_(net1483[14]),.decode_n14_VGRUN_2_(net1484[14]),.decode_n14_VGRUN_3_(net1485[14]),.decode_n15_VGRUN_0_(net1482[15]),.decode_n15_VGRUN_1_(net1483[15]),.decode_n15_VGRUN_2_(net1484[15]),.decode_n15_VGRUN_3_(net1485[15]));
	TSMC350nm_GateMuxSwcTile switch(.island_num(1), .direction(horizontal), .num(32));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect01d3 switch(.island_num(1), .direction(vertical), .num(16), .type(drain_select));
	TSMC350nm_FourTgate_ThickOx_FG_MEM switch(.island_num(1), .direction(vertical), .num(16), .type(prog_switch));
endmodule