module TOP(port1);


	/* Island 0 */
	TSMC350nm_C4 I__0 (.island_num(0), .row(0), .col(0), .matrix_row(12), .matrix_col(1), .OUTPUTcol_0(net268[0:12]));

 	/*Programming Mux */ 


	/* Island 1 */
	TSMC350nm_Ampdet_NoFG I__0 (.island_num(1), .row(0), .col(0), .matrix_row(12), .matrix_col(1), .VINcol_0(net268[0:12]), .OUTPUTcol_0(net280[0:12]));

 	/*Programming Mux */ 


	/* Island 2 */
	TSMC350nm_DelayBlock_3stage_new I__0 (.island_num(2), .row(0), .col(0), .matrix_row(12), .matrix_col(1), .VINcol_0(net280[0:12]));

 	/*Programming Mux */ 


	/* Island 3 */
	TSMC350nm_VMMWTA I__0 (.island_num(3), .row(0), .col(17), .matrix_row(9), .matrix_col(1), .matrix_row(9), .matrix_col(1));
	TSMC350nm_4x2_Indirect I__1 (.island_num(3), .row(0), .col(0), .matrix_row(9), .matrix_col(17));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(3), .direction(horizontal), .bits(6));
	TSMC350nm_IndirectSwitches switch(.island_num(3), .direction(horizontal), .num(18));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(3), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect01d3 switch(.island_num(3), .direction(vertical), .num(9), .type(drain_select));
	TSMC350nm_FourTgate_ThickOx_FG_MEM switch(.island_num(3), .direction(vertical), .num(9), .type(prog_switch));
endmodule