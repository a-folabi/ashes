module TOP(port1);


	/* Island 0 */
	TSMC350nm_TA2Cell_Weak I__0 (.island_num(0), .row(0), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net220[0]), .VD_P_1_row_0(net221[0]), .VIN1_PLUSrow_0(net297), .VIN1_MINUSrow_0(net30), .VIN2_PLUSrow_0(net30), .VIN2_MINUSrow_0(net71), .OUTPUT_0_row_0(net30), .OUTPUT_1_row_0(net30), .Vsel_0_row_0(net295), .Vsel_1_row_0(net296), .RUNrow_0(net323), .Vg_0_row_0(net293), .Vg_1_row_0(net294), .PROGrow_0(net322), .VTUNrow_0(net320), .VINJrow_0(net318), .GNDrow_0(net319), .VPWRrow_0(net321));
	TSMC350nm_TA2Cell_Weak I__1 (.island_num(0), .row(1), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net222[0]), .VD_P_1_row_0(net223[0]), .VIN1_PLUSrow_0(net30), .VIN1_MINUSrow_0(net71), .VIN2_PLUSrow_0(net71), .VIN2_MINUSrow_0(net299), .OUTPUT_0_row_0(net71), .OUTPUT_1_row_0(net299));
	TSMC350nm_TA2Cell_Weak I__2 (.island_num(0), .row(2), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net224[0]), .VD_P_1_row_0(net225[0]), .VIN1_PLUSrow_0(net71), .VIN1_MINUSrow_0(net72), .VIN2_PLUSrow_0(net72), .VIN2_MINUSrow_0(net113), .OUTPUT_0_row_0(net72), .OUTPUT_1_row_0(net72));
	TSMC350nm_TA2Cell_Weak I__3 (.island_num(0), .row(3), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net226[0]), .VD_P_1_row_0(net227[0]), .VIN1_PLUSrow_0(net72), .VIN1_MINUSrow_0(net113), .VIN2_PLUSrow_0(net113), .VIN2_MINUSrow_0(net300), .OUTPUT_0_row_0(net113), .OUTPUT_1_row_0(net300));
	TSMC350nm_TA2Cell_Weak I__4 (.island_num(0), .row(4), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net228[0]), .VD_P_1_row_0(net229[0]), .VIN1_PLUSrow_0(net113), .VIN1_MINUSrow_0(net114), .VIN2_PLUSrow_0(net114), .VIN2_MINUSrow_0(net155), .OUTPUT_0_row_0(net114), .OUTPUT_1_row_0(net114));
	TSMC350nm_TA2Cell_Weak I__5 (.island_num(0), .row(5), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net230[0]), .VD_P_1_row_0(net231[0]), .VIN1_PLUSrow_0(net114), .VIN1_MINUSrow_0(net155), .VIN2_PLUSrow_0(net155), .VIN2_MINUSrow_0(net301), .OUTPUT_0_row_0(net155), .OUTPUT_1_row_0(net301));
	TSMC350nm_TA2Cell_Weak I__6 (.island_num(0), .row(6), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net232[0]), .VD_P_1_row_0(net233[0]), .VIN1_PLUSrow_0(net155), .VIN1_MINUSrow_0(net156), .VIN2_PLUSrow_0(net156), .VIN2_MINUSrow_0(net195), .OUTPUT_0_row_0(net156), .OUTPUT_1_row_0(net156));
	TSMC350nm_TA2Cell_Weak I__7 (.island_num(0), .row(7), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net234[0]), .VD_P_1_row_0(net235[0]), .VIN1_PLUSrow_0(net156), .VIN1_MINUSrow_0(net195), .VIN2_PLUSrow_0(net195), .VIN2_MINUSrow_0(net302), .OUTPUT_0_row_0(net195), .OUTPUT_1_row_0(net302));
	TSMC350nm_TA2Cell_Weak I__8 (.island_num(0), .row(8), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net236[0]), .VD_P_1_row_0(net237[0]), .VIN1_PLUSrow_0(net195), .VIN1_MINUSrow_0(net196), .VIN2_PLUSrow_0(net196), .VIN2_MINUSrow_0(net298), .OUTPUT_0_row_0(net196), .OUTPUT_1_row_0(net196));
	TSMC350nm_TA2Cell_Weak I__9 (.island_num(0), .row(9), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net238[0]), .VD_P_1_row_0(net239[0]), .VIN1_PLUSrow_0(net196), .VIN1_MINUSrow_0(net298), .VIN2_PLUSrow_0(net298), .VIN2_MINUSrow_0(net303), .OUTPUT_0_row_0(net298), .OUTPUT_1_row_0(net303), .VINJ_brow_0(net317), .GND_brow_0(net316));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5), .decode_n0_IN_0_(net314), .decode_n2_IN_1_(net313), .decode_n2_IN_0_(net312), .decode_n4_IN_1_(net311), .decode_n4_IN_0_(net310), .decode_n0_ENABLE(net315));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select), .switch_n0_prog_drainrail(net309), .switch_n0_VINJ(net317), .switch_n0_GND(net316));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch), .switch_n0_PR_0_(net220[0]), .switch_n0_PR_1_(net221[0]), .switch_n0_PR_2_(net222[0]), .switch_n0_PR_3_(net223[0]), .switch_n1_PR_0_(net224[0]), .switch_n1_PR_1_(net225[0]), .switch_n1_PR_2_(net226[0]), .switch_n1_PR_3_(net227[0]), .switch_n2_PR_0_(net228[0]), .switch_n2_PR_1_(net229[0]), .switch_n2_PR_2_(net230[0]), .switch_n2_PR_3_(net231[0]), .switch_n3_PR_0_(net232[0]), .switch_n3_PR_1_(net233[0]), .switch_n3_PR_2_(net234[0]), .switch_n3_PR_3_(net235[0]), .switch_n4_PR_0_(net236[0]), .switch_n4_PR_1_(net237[0]), .switch_n4_PR_2_(net238[0]), .switch_n4_PR_3_(net239[0]), .switch_n0_VDD(net317), .switch_n0_GND(net316), .switch_n0_RUN(net323));
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(2), .decode_n0_ENABLE(net306), .decode_n0_VINJV(net318), .decode_n0_GNDV(net319), .decode_n0_n0_IN_1_(net308), .decode_n0_n0_IN_0_(net307));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(1));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(0), .direction(horizontal), .col(0), .RUN_IN_0_(net304), .RUN_IN_1_(net304), .GND_T(net319), .VINJ_T(net318), .CTRL_B_0_(net295), .CTRL_B_1_(net296), .Vg_0_(net293), .Vg_1_(net294), .PROG(net322), .RUN(net323), .Vgsel(net305));


	/* Frame */ 
	tile_analog_frame cab_frame(.pin_layer(METAL3), .W_w_Vin(net297), .E_e_Vout(net298), .E_e_Vout_Buf_0_(net299), .E_e_Vout_Buf_1_(net300), .E_e_Vout_Buf_2_(net301), .E_e_Vout_Buf_3_(net302), .E_e_Vout_Buf_4_(net303), .N_n_Prog(net322), .N_n_Run(net323), .N_n_VGRUN(net304), .N_n_VGPROG(net305), .N_n_VTUN(net320), .N_n_AVDD(net321), .N_n_gnd(net319), .S_s_gnd(net316), .N_n_vinj(net318), .S_s_vinj(net317), .S_s_Drainline_Prog(net309), .N_n_GateEnable(net306), .W_w_GateB_0_(net307), .W_w_GateB_1_(net308), .W_w_DrainEnable(net315), .W_w_DrainB_0_(net310), .W_w_DrainB_1_(net311), .W_w_DrainB_2_(net312), .W_w_DrainB_3_(net313), .W_w_DrainB_4_(net314));
 endmodule