module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(7), .GND_b_1_row_4(net2359[0:7]), .Vs_b_0_row_4(net124[0:7]), .Vs_b_1_row_4(net125[0:7]), .VINJ_b_1_row_4(net2366[0:7]), .Vsel_b_0_row_4(net2324[0:7]), .Vsel_b_1_row_4(net2325[0:7]), .Vg_b_0_row_4(net2338[0:7]), .Vg_b_1_row_4(net2339[0:7]), .VTUN_brow_4(net2352[0:7]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(17), .matrix_row(5), .matrix_col(9), .GND_b_1_row_4(net2402[0:9]), .Vs_b_0_row_4(net325[0:9]), .Vs_b_1_row_4(net326[0:9]), .VINJ_b_1_row_4(net2401[0:9]), .Vsel_b_0_row_4(net2403[0:9]), .Vsel_b_1_row_4(net2405[0:9]), .Vg_b_0_row_4(net344[0:9]), .Vg_b_1_row_4(net345[0:9]), .VTUN_brow_4(net2400[0:9]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(26), .matrix_row(5), .matrix_col(1), .Prog_brow_4(net2574[0:1]), .VDD_brow_4(net2573[0:1]), .GND_brow_4(net2402[8:9]));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2379[0:1]), .Vsel_b_0_row_4(net2382[0:1]), .Vsel_b_1_row_4(net2383[0:1]), .Vg_b_0_row_4(net2384[0:1]), .Vg_b_1_row_4(net2385[0:1]), .VTUN_brow_4(net2380[0:1]), .GND_b_1_row_4(net2381[0:1]));
	S_BLOCK_BUFFER I__4 (.island_num(0), .row(0), .col(8), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__5 (.island_num(0), .row(0), .col(9), .matrix_row(4), .matrix_col(1));
	S_BLOCK_CONN_PINS I__6 (.island_num(0), .row(4), .col(9), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__7 (.island_num(0), .row(0), .col(10), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__8 (.island_num(0), .row(3), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__9 (.island_num(0), .row(4), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__10 (.island_num(0), .row(0), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_CONN_PINS I__11 (.island_num(0), .row(2), .col(11), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__12 (.island_num(0), .row(3), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__13 (.island_num(0), .row(0), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_CONN_PINS I__14 (.island_num(0), .row(1), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__15 (.island_num(0), .row(2), .col(12), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__16 (.island_num(0), .row(0), .col(13), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__17 (.island_num(0), .row(1), .col(13), .matrix_row(4), .matrix_col(1));
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2386[0:1]), .Vsel_b_0_row_4(net2389[0:1]), .Vsel_b_1_row_4(net2390[0:1]), .Vg_b_0_row_4(net2391[0:1]), .Vg_b_1_row_4(net2392[0:1]), .VTUN_brow_4(net2387[0:1]), .GND_b_1_row_4(net2388[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2393[0:1]), .Vsel_b_0_row_4(net2396[0:1]), .Vsel_b_1_row_4(net2397[0:1]), .Vg_b_0_row_4(net2398[0:1]), .Vg_b_1_row_4(net2399[0:1]), .VTUN_brow_4(net2394[0:1]), .GND_b_1_row_4(net2395[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(6), .decode_n0_VINJ_b_0_(net2401[8]), .decode_n0_VINJ_b_1_(net2401[8]), .decode_n1_VINJ_b_0_(net2401[8]), .decode_n1_VINJ_b_1_(net2401[8]), .decode_n2_VINJ_b_0_(net2401[8]), .decode_n2_VINJ_b_1_(net2401[8]), .decode_n3_VINJ_b_0_(net2401[8]), .decode_n3_VINJ_b_1_(net2401[8]), .decode_n4_VINJ_b_1_(net2468), .decode_n5_VINJ_b_0_(net2470), .decode_n5_VINJ_b_1_(net2472), .decode_n6_VINJ_b_0_(net2474), .decode_n6_VINJ_b_1_(net2476), .decode_n7_VINJ_b_0_(net2478), .decode_n7_VINJ_b_1_(net2480), .decode_n8_VINJ_b_0_(net2482), .decode_n8_VINJ_b_1_(net2484), .decode_n9_VINJ_b_0_(net2486), .decode_n9_VINJ_b_1_(net2488), .decode_n0_GND_b_0_(net2402[8]), .decode_n0_GND_b_1_(net2402[8]), .decode_n1_GND_b_0_(net2402[8]), .decode_n1_GND_b_1_(net2402[8]), .decode_n2_GND_b_0_(net2402[8]), .decode_n2_GND_b_1_(net2402[8]), .decode_n3_GND_b_0_(net2402[8]), .decode_n3_GND_b_1_(net2402[8]), .decode_n4_GND_b_1_(net2469), .decode_n5_GND_b_0_(net2471), .decode_n5_GND_b_1_(net2473), .decode_n6_GND_b_0_(net2475), .decode_n6_GND_b_1_(net2477), .decode_n7_GND_b_0_(net2479), .decode_n7_GND_b_1_(net2481), .decode_n8_GND_b_0_(net2483), .decode_n8_GND_b_1_(net2485), .decode_n9_GND_b_0_(net2487), .decode_n9_GND_b_1_(net2489));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(26), .switch_n0_RUN_IN_0_(net2575[0]), .switch_n0_RUN_IN_1_(net2575[0]), .switch_n1_RUN_IN_0_(net2575[0]), .switch_n1_RUN_IN_1_(net2575[0]), .switch_n2_RUN_IN_0_(net2575[0]), .switch_n2_RUN_IN_1_(net2575[0]), .switch_n3_RUN_IN_0_(net2575[0]), .switch_n3_RUN_IN_1_(net2575[0]), .switch_n4_RUN_IN_0_(net2575[0]), .switch_n4_RUN_IN_1_(net2575[0]), .switch_n5_RUN_IN_0_(net2575[0]), .switch_n5_RUN_IN_1_(net2575[0]), .switch_n6_RUN_IN_0_(net2575[0]), .switch_n6_RUN_IN_1_(net2575[0]), .switch_n7_RUN_IN_0_(net2575[0]), .switch_n7_RUN_IN_1_(net2575[0]), .switch_n14_RUN_IN_0_(net2575[0]), .switch_n14_RUN_IN_1_(net2575[0]), .switch_n16_RUN_IN_0_(net2575[0]), .switch_n16_RUN_IN_1_(net2575[0]), .switch_n17_RUN_IN_0_(net2575[0]), .switch_n17_RUN_IN_1_(net2575[0]), .switch_n18_RUN_IN_0_(net2575[0]), .switch_n18_RUN_IN_1_(net2575[0]), .switch_n19_RUN_IN_0_(net2575[0]), .switch_n19_RUN_IN_1_(net2575[0]), .switch_n20_RUN_IN_0_(net2575[0]), .switch_n20_RUN_IN_1_(net2575[0]), .switch_n21_RUN_IN_0_(net2575[0]), .switch_n21_RUN_IN_1_(net2575[0]), .switch_n22_RUN_IN_0_(net2575[0]), .switch_n22_RUN_IN_1_(net2575[0]), .switch_n23_RUN_IN_0_(net2575[0]), .switch_n23_RUN_IN_1_(net2575[0]), .switch_n24_RUN_IN_0_(net2575[0]), .switch_n24_RUN_IN_1_(net2575[0]), .switch_n25_RUN_IN_0_(net2575[0]), .switch_n25_RUN_IN_1_(net2575[0]), .switch_n14_GND_T(net2469), .switch_n16_GND_T(net2471), .switch_n17_GND_T(net2473), .switch_n18_GND_T(net2475), .switch_n19_GND_T(net2477), .switch_n20_GND_T(net2479), .switch_n21_GND_T(net2481), .switch_n22_GND_T(net2483), .switch_n23_GND_T(net2485), .switch_n24_GND_T(net2487), .switch_n25_GND_T(net2489), .switch_n14_VINJ_T(net2468), .switch_n16_VINJ_T(net2470), .switch_n17_VINJ_T(net2472), .switch_n18_VINJ_T(net2474), .switch_n19_VINJ_T(net2476), .switch_n20_VINJ_T(net2478), .switch_n21_VINJ_T(net2480), .switch_n22_VINJ_T(net2482), .switch_n23_VINJ_T(net2484), .switch_n24_VINJ_T(net2486), .switch_n25_VINJ_T(net2488));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch));
	none switch_ind(.island_num(0), .direction(horizontal), .col(8));
	none switch_ind(.island_num(0), .direction(horizontal), .col(9));
	none switch_ind(.island_num(0), .direction(horizontal), .col(10));
	none switch_ind(.island_num(0), .direction(horizontal), .col(11));
	none switch_ind(.island_num(0), .direction(horizontal), .col(12));
	none switch_ind(.island_num(0), .direction(horizontal), .col(13));
	none switch_ind(.island_num(0), .direction(horizontal), .col(15));


	/* Island 1 */
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__0 (.island_num(1), .row(0), .col(0), .matrix_row(1), .matrix_col(8));
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(7), .matrix_col(8), .GND_b_0_row_6(net1353[0:8]), .GND_b_1_row_6(net1354[0:8]), .Vs_b_0_row_6(net1363[0:8]), .Vs_b_1_row_6(net1364[0:8]), .VINJ_b_0_row_6(net1367[0:8]), .VINJ_b_1_row_6(net1368[0:8]), .Vsel_b_0_row_6(net1371[0:8]), .Vsel_b_1_row_6(net1372[0:8]), .Vg_b_0_row_6(net1375[0:8]), .Vg_b_1_row_6(net1376[0:8]), .VTUN_brow_6(net1379[0:8]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(8), .matrix_row(6), .matrix_col(10));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(7), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2226), .P_1_row_0(net2227), .A_0_row_0(net2228), .A_1_row_0(net2229), .A_2_row_0(net2230), .A_3_row_0(net2231));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2238), .P_1_row_0(net2239), .A_0_row_0(net2240), .A_1_row_0(net2241), .A_2_row_0(net2242), .A_3_row_0(net2243));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2256), .P_1_row_0(net2257), .A_0_row_0(net2258), .A_1_row_0(net2259), .A_2_row_0(net2260), .A_3_row_0(net2261));
	TSMC350nm_4TGate_ST_BMatrix_NoSwitch I__8 (.island_num(1), .row(3), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2274), .P_1_row_0(net2275), .P_2_row_0(net2276), .P_3_row_0(net2277), .A_0_row_0(net2278), .A_1_row_0(net2279), .A_2_row_0(net2280), .A_3_row_0(net2281));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2293), .P_1_row_0(net2294), .P_2_row_0(net2295), .P_3_row_0(net2296), .A_0_row_0(net2297), .A_1_row_0(net2298));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net2308), .A_1_row_0(net2309), .A_2_row_0(net2310), .A_3_row_0(net2311));
	TSMC350nm_4TGate_ST_BMatrix I__11 (.island_num(1), .row(6), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net2315), .A_1_row_0(net2316), .A_2_row_0(net2317), .A_3_row_0(net2318));
	TSMC350nm_4TGate_ST_BMatrix I__12 (.island_num(1), .row(7), .col(18), .matrix_row(1), .matrix_col(1), .Prog_brow_0(net2574[0]), .VDD_brow_0(net2573[0]), .GND_brow_0(net2402[8]));
	TSMC350nm_OutMtrx_IndrctSwcs I__13 (.island_num(1), .row(9), .col(8), .matrix_row(1), .matrix_col(10), .Vgrun_rcol_9(net2575[0:1]), .AVDD_rcol_9(net2569[0:1]), .run_rcol_9(net2571[0:1]), .prog_rcol_9(net2570[0:1]));
	TSMC350nm_4x2_Indirect I__14 (.island_num(1), .row(10), .col(8), .matrix_row(2), .matrix_col(10), .Vd_Rl_0_col_0(net2063[0:2]), .Vd_Rl_1_col_0(net2064[0:2]), .Vd_Rl_2_col_0(net2065[0:2]), .Vd_Rl_3_col_0(net2066[0:2]), .Vd_Pl_0_col_0(net2067[0:2]), .Vd_Pl_1_col_0(net2068[0:2]), .Vd_Pl_2_col_0(net2069[0:2]), .Vd_Pl_3_col_0(net2070[0:2]));
	TSMC350nm_4TGate_ST_BMatrix I__15 (.island_num(1), .row(10), .col(18), .matrix_row(2), .matrix_col(1), .Prog_brow_1(net2574[0:1]), .VDD_brow_1(net2573[0:1]), .GND_brow_1(net2402[8:9]));
	TSMC350nm_TA2Cell_Weak cab_device_16 (.island_num(1), .row(2), .col(19), .VD_P_0_(net2226), .VD_P_1_(net2227), .VIN1_PLUS(net2228), .VIN1_MINUS(net2229), .VIN2_PLUS(net2230), .VIN2_MINUS(net2231), .OUTPUT_0_(net2232[0]), .OUTPUT_1_(net2233[0]), .Vsel_0_(net2302), .Vsel_1_(net2303), .RUN(net2234), .Vg_0_(net2304), .Vg_1_(net2305), .PROG(net2574[0]), .VTUN(net2235), .VINJ(net2236), .GND(net2237), .VPWR(net2569[0]), .Vsel_b_0_(net2246), .Vsel_b_1_(net2247), .RUN_b(net2248), .Vg_b_0_(net2249), .Vg_b_1_(net2250), .PROG_b(net2251), .VTUN_b(net2252), .VINJ_b(net2253), .GND_b(net2254), .VPWR_b(net2255));
	TSMC350nm_TA2Cell_Weak cab_device_17 (.island_num(1), .row(3), .col(19), .VD_P_0_(net2238), .VD_P_1_(net2239), .VIN1_PLUS(net2240), .VIN1_MINUS(net2241), .VIN2_PLUS(net2242), .VIN2_MINUS(net2243), .OUTPUT_0_(net2244[0]), .OUTPUT_1_(net2245[0]), .Vsel_0_(net2246), .Vsel_1_(net2247), .RUN(net2248), .Vg_0_(net2249), .Vg_1_(net2250), .PROG(net2251), .VTUN(net2252), .VINJ(net2253), .GND(net2254), .VPWR(net2255), .Vsel_b_0_(net2264), .Vsel_b_1_(net2265), .RUN_b(net2266), .Vg_b_0_(net2267), .Vg_b_1_(net2268), .PROG_b(net2269), .VTUN_b(net2270), .VINJ_b(net2271), .GND_b(net2272), .VPWR_b(net2273));
	TSMC350nm_TA2Cell_Strong cab_device_18 (.island_num(1), .row(4), .col(19), .VD_P_0_(net2256), .VD_P_1_(net2257), .VIN1_PLUS(net2258), .VIN1_MINUS(net2259), .VIN2_PLUS(net2260), .VIN2_MINUS(net2261), .OUTPUT_0_(net2262[0]), .OUTPUT_1_(net2263[0]), .Vsel_0_(net2264), .Vsel_1_(net2265), .RUN(net2266), .Vg_0_(net2267), .Vg_1_(net2268), .PROG(net2269), .VTUN(net2270), .VINJ(net2271), .GND(net2272), .VPWR(net2273), .Vg_b_0_(net2289), .PROG_b(net2292), .VTUN_b(net2290), .VINJ_b(net2288), .GND_b(net2291));
	TSMC350nm_4WTA_IndirectProg cab_device_19 (.island_num(1), .row(5), .col(19), .VD_P_0_(net2274), .VD_P_1_(net2275), .VD_P_2_(net2276), .VD_P_3_(net2277), .Iin_0_(net2278), .Iin_1_(net2279), .Iin_2_(net2280), .Iin_3_(net2281), .Vout_0_(net2282[0]), .Vout_1_(net2283[0]), .Vout_2_(net2284[0]), .Vout_3_(net2285[0]), .Vmid(net2286[0]), .Vbias(net2287[0]), .Vsel(net2302), .Vs(net2569[0]), .VINJ(net2288), .Vg(net2289), .VTUN(net2290), .GND(net2291), .PROG(net2292), .VINJ_b(net2301), .VTUN_b(net2307), .GND_b(net2306));
	TSMC350nm_Cap_Bank cab_device_20 (.island_num(1), .row(6), .col(19), .VD_P_0_(net2293), .VD_P_1_(net2294), .VD_P_2_(net2295), .VD_P_3_(net2296), .VIN_0_(net2297), .VIN_1_(net2298), .OUT_0_(net2299[0]), .OUT_1_(net2300[0]), .VINJ(net2301), .Vsel_0_(net2302), .Vsel_1_(net2303), .Vg_0_(net2304), .Vg_1_(net2305), .GND(net2306), .VTUN(net2307), .GND_b(net2314));
	TSMC350nm_NandPfets cab_device_21 (.island_num(1), .row(7), .col(19), .GATE_N(net2308), .SOURCE_N(net2309), .GATE_P(net2310), .SOURCE_P(net2311), .DRAIN_N(net2312[0]), .DRAIN_P(net2313[0]), .VPWR(net2569[0]), .GND(net2314), .VPWR_b(net2322), .GND_b(net2323));
	TSMC350nm_TGate_2nMirror cab_device_22 (.island_num(1), .row(8), .col(19), .IN_CM_0_(net2315), .IN_CM_1_(net2316), .SelN(net2317), .IN_TG(net2318), .OUT_CM_0_(net2319[0]), .OUT_CM_1_(net2320[0]), .OUT_TG(net2321[0]), .VPWR(net2322), .GND(net2323));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(1), .direction(vertical), .num(12), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(12), .type(prog_switch), .switch_n8_PR_0_(net2554[0]), .switch_n8_PR_1_(net2558[0]), .switch_n8_PR_2_(net2562[0]), .switch_n8_PR_3_(net2566[0]), .switch_n8_In_0_(net2553[0]), .switch_n8_In_1_(net2557[0]), .switch_n8_In_2_(net2561[0]), .switch_n8_In_3_(net2565[0]));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(20), .switch_n0_Input_0_(net2573[0]), .switch_n0_Input_1_(net2359[0]), .switch_n1_Input_0_(net124[1]), .switch_n1_Input_1_(net125[1]), .switch_n2_Input_0_(net124[2]), .switch_n2_Input_1_(net125[2]), .switch_n3_Input_0_(net124[3]), .switch_n3_Input_1_(net125[3]), .switch_n4_Input_0_(net325[0]), .switch_n4_Input_1_(net326[0]), .switch_n5_Input_0_(net325[1]), .switch_n5_Input_1_(net326[1]), .switch_n6_Input_0_(net325[2]), .switch_n6_Input_1_(net326[2]), .switch_n7_Input_0_(net325[3]), .switch_n7_Input_1_(net326[3]), .switch_n8_Input_0_(net2552[0]), .switch_n8_Input_1_(net2232[0]), .switch_n9_Input_0_(net2233[0]), .switch_n9_Input_1_(net2244[0]), .switch_n10_Input_0_(net2245[0]), .switch_n10_Input_1_(net2262[0]), .switch_n11_Input_0_(net2263[0]), .switch_n11_Input_1_(net2282[0]), .switch_n12_Input_0_(net2283[0]), .switch_n12_Input_1_(net2284[0]), .switch_n13_Input_0_(net2285[0]), .switch_n13_Input_1_(net2286[0]), .switch_n14_Input_0_(net2287[0]), .switch_n14_Input_1_(net2299[0]), .switch_n15_Input_0_(net2300[0]), .switch_n15_Input_1_(net2312[0]), .switch_n16_Input_0_(net2313[0]), .switch_n16_Input_1_(net2319[0]), .switch_n17_Input_0_(net2320[0]), .switch_n17_Input_1_(net2321[0]), .switch_n0_GND(net2359[0]), .switch_n1_GND(net2359[1]), .switch_n2_GND(net2359[2]), .switch_n3_GND(net2359[3]), .switch_n4_GND(net2359[4]), .switch_n5_GND(net2359[5]), .switch_n6_GND(net2359[6]), .switch_n7_GND(net2381[0]), .switch_n8_GND(net2388[0]), .switch_n9_GND(net2395[0]), .switch_n10_GND(net2402[0]), .switch_n11_GND(net2402[1]), .switch_n12_GND(net2402[2]), .switch_n13_GND(net2402[3]), .switch_n14_GND(net2402[4]), .switch_n15_GND(net2402[5]), .switch_n16_GND(net2402[6]), .switch_n17_GND(net2402[7]), .switch_n0_Vsel_0_(net2324[0]), .switch_n0_Vsel_1_(net2325[0]), .switch_n1_Vsel_0_(net2324[1]), .switch_n1_Vsel_1_(net2325[1]), .switch_n2_Vsel_0_(net2324[2]), .switch_n2_Vsel_1_(net2325[2]), .switch_n3_Vsel_0_(net2324[3]), .switch_n3_Vsel_1_(net2325[3]), .switch_n4_Vsel_0_(net2324[4]), .switch_n4_Vsel_1_(net2325[4]), .switch_n5_Vsel_0_(net2324[5]), .switch_n5_Vsel_1_(net2325[5]), .switch_n6_Vsel_0_(net2324[6]), .switch_n6_Vsel_1_(net2325[6]), .switch_n7_Vsel_0_(net2383[0]), .switch_n7_Vsel_1_(net2382[0]), .switch_n8_Vsel_0_(net2390[0]), .switch_n8_Vsel_1_(net2389[0]), .switch_n9_Vsel_0_(net2397[0]), .switch_n9_Vsel_1_(net2396[0]), .switch_n10_Vsel_0_(net2403[0]), .switch_n10_Vsel_1_(net2405[0]), .switch_n11_Vsel_0_(net2403[1]), .switch_n11_Vsel_1_(net2405[1]), .switch_n12_Vsel_0_(net2403[2]), .switch_n12_Vsel_1_(net2405[2]), .switch_n13_Vsel_0_(net2403[3]), .switch_n13_Vsel_1_(net2405[3]), .switch_n14_Vsel_0_(net2403[4]), .switch_n14_Vsel_1_(net2405[4]), .switch_n15_Vsel_0_(net2403[5]), .switch_n15_Vsel_1_(net2405[5]), .switch_n16_Vsel_0_(net2403[6]), .switch_n16_Vsel_1_(net2405[6]), .switch_n17_Vsel_0_(net2403[7]), .switch_n17_Vsel_1_(net2405[7]), .switch_n0_Vg_global_0_(net2338[0]), .switch_n0_Vg_global_1_(net2339[0]), .switch_n1_Vg_global_0_(net2338[1]), .switch_n1_Vg_global_1_(net2339[1]), .switch_n2_Vg_global_0_(net2338[2]), .switch_n2_Vg_global_1_(net2339[2]), .switch_n3_Vg_global_0_(net2338[3]), .switch_n3_Vg_global_1_(net2339[3]), .switch_n4_Vg_global_0_(net2338[4]), .switch_n4_Vg_global_1_(net2339[4]), .switch_n5_Vg_global_0_(net2338[5]), .switch_n5_Vg_global_1_(net2339[5]), .switch_n6_Vg_global_0_(net2338[6]), .switch_n6_Vg_global_1_(net2339[6]), .switch_n7_Vg_global_0_(net2385[0]), .switch_n7_Vg_global_1_(net2384[0]), .switch_n8_Vg_global_0_(net2392[0]), .switch_n8_Vg_global_1_(net2391[0]), .switch_n9_Vg_global_0_(net2399[0]), .switch_n9_Vg_global_1_(net2398[0]), .switch_n10_Vg_global_0_(net344[0]), .switch_n10_Vg_global_1_(net345[0]), .switch_n11_Vg_global_0_(net344[1]), .switch_n11_Vg_global_1_(net345[1]), .switch_n12_Vg_global_0_(net344[2]), .switch_n12_Vg_global_1_(net345[2]), .switch_n13_Vg_global_0_(net344[3]), .switch_n13_Vg_global_1_(net345[3]), .switch_n14_Vg_global_0_(net344[4]), .switch_n14_Vg_global_1_(net345[4]), .switch_n15_Vg_global_0_(net344[5]), .switch_n15_Vg_global_1_(net345[5]), .switch_n16_Vg_global_0_(net344[6]), .switch_n16_Vg_global_1_(net345[6]), .switch_n17_Vg_global_0_(net344[7]), .switch_n17_Vg_global_1_(net345[7]), .switch_n0_VTUN(net2352[0]), .switch_n1_VTUN(net2352[1]), .switch_n2_VTUN(net2352[2]), .switch_n3_VTUN(net2352[3]), .switch_n4_VTUN(net2352[4]), .switch_n5_VTUN(net2352[5]), .switch_n6_VTUN(net2352[6]), .switch_n7_VTUN(net2380[0]), .switch_n8_VTUN(net2387[0]), .switch_n9_VTUN(net2394[0]), .switch_n10_VTUN(net2400[0]), .switch_n11_VTUN(net2400[1]), .switch_n12_VTUN(net2400[2]), .switch_n13_VTUN(net2400[3]), .switch_n14_VTUN(net2400[4]), .switch_n15_VTUN(net2400[5]), .switch_n16_VTUN(net2400[6]), .switch_n17_VTUN(net2400[7]), .switch_n0_VINJ(net2366[0]), .switch_n1_VINJ(net2366[1]), .switch_n2_VINJ(net2366[2]), .switch_n3_VINJ(net2366[3]), .switch_n4_VINJ(net2366[4]), .switch_n5_VINJ(net2366[5]), .switch_n6_VINJ(net2366[6]), .switch_n7_VINJ(net2379[0]), .switch_n8_VINJ(net2386[0]), .switch_n9_VINJ(net2393[0]), .switch_n10_VINJ(net2401[0]), .switch_n11_VINJ(net2401[1]), .switch_n12_VINJ(net2401[2]), .switch_n13_VINJ(net2401[3]), .switch_n14_VINJ(net2401[4]), .switch_n15_VINJ(net2401[5]), .switch_n16_VINJ(net2401[6]), .switch_n17_VINJ(net2401[7]), .switch_n0_Vgrun_r(net2575[0]), .switch_n0_AVDD_r(net2569[0]), .switch_n0_run_r(net2571[0]), .switch_n0_prog_r(net2570[0]));
	none switch_ind(.island_num(1), .direction(horizontal), .col(18));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(19), .VPWR_0_(net2573[0]), .VPWR_1_(net2573[0]), .RUN_IN_0_(net2575[0]), .RUN_IN_1_(net2575[0]), .GND_T(net2402[8]), .VTUN_T(net2400[8]), .decode_0_(net2403[8]), .decode_1_(net2405[8]), .VINJ_T(net2401[8]), .GND(net2237), .CTRL_B_0_(net2302), .CTRL_B_1_(net2303), .run_r(net2234), .prog_r(net2574[0]), .Vg_0_(net2304), .Vg_1_(net2305), .VTUN(net2235), .VINJ(net2236), .VDD_1_(net2569[0]), .PROG(net2570[0]), .RUN(net2571[0]));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net1363[0:6]), .out_1_row_0(net1364[0:6]), .VINJ_0_row_0(net1367[0:6]), .VINJ_1_row_0(net1368[0:6]), .Vsel_0_row_0(net1371[0:6]), .Vsel_1_row_0(net1372[0:6]), .Vg_0_row_0(net1375[0:6]), .Vg_1_row_0(net1376[0:6]), .GNDrow_0(net1353[0:6]), .VTUNrow_0(net1379[0:6]), .Dcol_0(net124[6:7]), .CLKcol_0(net125[6:7]), .Qcol_5(net125[6:7]), .comcol_0(net2552[0:1]), .VDDcol_0(net2569[0:1]), .Vd_Pcol_0(net2566[0:1]), .Vd_in_0_col_0(net2553[0:1]), .Vd_in_1_col_0(net2557[0:1]), .Vd_in_2_col_0(net2561[0:1]), .Vd_in_3_col_0(net2565[0:1]), .Vd_in_4_col_0(net2554[0:1]), .Vd_in_5_col_0(net2558[0:1]), .Vd_in_6_col_0(net2562[0:1]), .Vd_in_7_col_0(net2566[0:1]), .Vd_o_0_col_5(net2063[0:1]), .Vd_o_1_col_5(net2064[0:1]), .Vd_o_2_col_5(net2065[0:1]), .Vd_o_3_col_5(net2066[0:1]), .Vd_o_4_col_5(net2067[0:1]), .Vd_o_5_col_5(net2068[0:1]), .Vd_o_6_col_5(net2069[0:1]), .Vd_o_7_col_5(net2070[0:1]));

 	/*Programming Mux */ 


	/* Frame */ 
	tile_analog_frame cab_frame(.pin_layer(METAL3));
 endmodule