VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER routingPitch REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.01 ;
LAYER POLY1
  TYPE MASTERSLICE ;
END POLY1

LAYER CONT
  TYPE CUT ;
  SPACING 0.4 ;
END CONT

LAYER METAL1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.5 ;
  SPACING 0.45 ;
  PROPERTY routingPitch 1.25 ;
END METAL1

LAYER VIA12
  TYPE CUT ;
  SPACING 0.45 ;
END VIA12

LAYER METAL2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.4 ;
END METAL2

LAYER VIA23
  TYPE CUT ;
  SPACING 0.45 ;
END VIA23

LAYER METAL3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.25 ;
END METAL3

LAYER VIA34
  TYPE CUT ;
  SPACING 0.45 ;
END VIA34

LAYER METAL4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.6 ;
  PROPERTY routingPitch 1.4 ;
END METAL4

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIARULE M4_M3 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL4 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1

VIARULE M1_POLY1 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 1 ;
END M1_POLY1

VIA M1_POLY1
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER POLY1 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.35 -0.35 0.35 0.35 ;
END M1_POLY1

VIA M2_M1
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL2 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M2_M1

VIA M3_M2
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL3 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL2 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M3_M2

VIA M4_M3
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL3 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M4_M3


MACRO cab1
  PIN n_gateEN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 13.3 564.59 14.7 567.39 ;
    END
  END n_gateEN
  PIN n_programdrain
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 27.3 564.59 28.7 567.39 ;
    END
  END n_programdrain
  PIN n_rundrain
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 41.3 564.59 42.7 567.39 ;
    END
  END n_rundrain
  PIN n_cew0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 55.3 564.59 56.7 567.39 ;
    END
  END n_cew0
  PIN n_cew1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 69.3 564.59 70.7 567.39 ;
    END
  END n_cew1
  PIN n_cew2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 83.3 564.59 84.7 567.39 ;
    END
  END n_cew2
  PIN n_cew3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.3 564.59 98.7 567.39 ;
    END
  END n_cew3
  PIN n_vtun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 111.3 564.59 112.7 567.39 ;
    END
  END n_vtun
  PIN n_vinj<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 125.3 564.59 126.7 567.39 ;
    END
  END n_vinj<0>
  PIN n_vinj<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 139.3 564.59 140.7 567.39 ;
    END
  END n_vinj<1>
  PIN n_vinj<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 153.3 564.59 154.7 567.39 ;
    END
  END n_vinj<2>
  PIN n_gnd<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 167.3 564.59 168.7 567.39 ;
    END
  END n_gnd<0>
  PIN n_gnd<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 181.3 564.59 182.7 567.39 ;
    END
  END n_gnd<1>
  PIN n_gnd<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 195.3 564.59 196.7 567.39 ;
    END
  END n_gnd<2>
  PIN n_avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 209.3 564.59 210.7 567.39 ;
    END
  END n_avdd
  PIN n_s0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 223.3 564.59 224.7 567.39 ;
    END
  END n_s0
  PIN n_s1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 237.3 564.59 238.7 567.39 ;
    END
  END n_s1
  PIN n_s2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 251.3 564.59 252.7 567.39 ;
    END
  END n_s2
  PIN n_s3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 265.3 564.59 266.7 567.39 ;
    END
  END n_s3
  PIN n_s4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 279.3 564.59 280.7 567.39 ;
    END
  END n_s4
  PIN n_s5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 293.3 564.59 294.7 567.39 ;
    END
  END n_s5
  PIN n_s6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 307.3 564.59 308.7 567.39 ;
    END
  END n_s6
  PIN n_s7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 321.3 564.59 322.7 567.39 ;
    END
  END n_s7
  PIN n_s8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 335.3 564.59 336.7 567.39 ;
    END
  END n_s8
  PIN n_s9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 349.3 564.59 350.7 567.39 ;
    END
  END n_s9
  PIN n_s10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 363.3 564.59 364.7 567.39 ;
    END
  END n_s10
  PIN n_s11
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 377.3 564.59 378.7 567.39 ;
    END
  END n_s11
  PIN n_prog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 391.3 564.59 392.7 567.39 ;
    END
  END n_prog
  PIN n_run
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 405.3 564.59 406.7 567.39 ;
    END
  END n_run
  PIN n_vgsel
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 419.3 564.59 420.7 567.39 ;
    END
  END n_vgsel
  PIN e_cns0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 551.99 875.45 553.39 ;
    END
  END e_cns0
  PIN e_cns1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 537.99 875.45 539.39 ;
    END
  END e_cns1
  PIN e_cns2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 523.99 875.45 525.39 ;
    END
  END e_cns2
  PIN e_cns3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 509.99 875.45 511.39 ;
    END
  END e_cns3
  PIN e_vgrun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 495.99 875.45 497.39 ;
    END
  END e_vgrun
  PIN e_vtun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 481.99 875.45 483.39 ;
    END
  END e_vtun
  PIN e_vinj
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 467.99 875.45 469.39 ;
    END
  END e_vinj
  PIN e_gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 453.99 875.45 455.39 ;
    END
  END e_gnd
  PIN e_avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 439.99 875.45 441.39 ;
    END
  END e_avdd
  PIN e_drainbit3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 425.99 875.45 427.39 ;
    END
  END e_drainbit3
  PIN e_drainbit2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 411.99 875.45 413.39 ;
    END
  END e_drainbit2
  PIN e_drainbit1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 397.99 875.45 399.39 ;
    END
  END e_drainbit1
  PIN e_drainbit0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 383.99 875.45 385.39 ;
    END
  END e_drainbit0
  PIN e_s0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 369.99 875.45 371.39 ;
    END
  END e_s0
  PIN e_s1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 355.99 875.45 357.39 ;
    END
  END e_s1
  PIN e_s2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 341.99 875.45 343.39 ;
    END
  END e_s2
  PIN e_s3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 327.99 875.45 329.39 ;
    END
  END e_s3
  PIN e_s4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 313.99 875.45 315.39 ;
    END
  END e_s4
  PIN e_s5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 299.99 875.45 301.39 ;
    END
  END e_s5
  PIN e_s6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 285.99 875.45 287.39 ;
    END
  END e_s6
  PIN e_s7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 271.99 875.45 273.39 ;
    END
  END e_s7
  PIN e_s8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 257.99 875.45 259.39 ;
    END
  END e_s8
  PIN e_s9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 243.99 875.45 245.39 ;
    END
  END e_s9
  PIN e_s10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 229.99 875.45 231.39 ;
    END
  END e_s10
  PIN e_s11
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 215.99 875.45 217.39 ;
    END
  END e_s11
  PIN e_drainbit9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 201.99 875.45 203.39 ;
    END
  END e_drainbit9
  PIN e_drainbit8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 187.99 875.45 189.39 ;
    END
  END e_drainbit8
  PIN e_drainbit7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 173.99 875.45 175.39 ;
    END
  END e_drainbit7
  PIN e_drainbit6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 159.99 875.45 161.39 ;
    END
  END e_drainbit6
  PIN e_drainbit5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 145.99 875.45 147.39 ;
    END
  END e_drainbit5
  PIN e_drainbit4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 131.99 875.45 133.39 ;
    END
  END e_drainbit4
  PIN e_drainEN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 117.99 875.45 119.39 ;
    END
  END e_drainEN
  PIN s_gateEN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 13.3 0.0 14.7 2.8 ;
    END
  END s_gateEN
  PIN s_programdrain
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 27.3 0.0 28.7 2.8 ;
    END
  END s_programdrain
  PIN s_rundrain
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 41.3 0.0 42.7 2.8 ;
    END
  END s_rundrain
  PIN s_cew0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 55.3 0.0 56.7 2.8 ;
    END
  END s_cew0
  PIN s_cew1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 69.3 0.0 70.7 2.8 ;
    END
  END s_cew1
  PIN s_cew2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 83.3 0.0 84.7 2.8 ;
    END
  END s_cew2
  PIN s_cew3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.3 0.0 98.7 2.8 ;
    END
  END s_cew3
  PIN s_vtun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 111.3 0.0 112.7 2.8 ;
    END
  END s_vtun
  PIN s_vinj<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 125.3 0.0 126.7 2.8 ;
    END
  END s_vinj<0>
  PIN s_vinj<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 139.3 0.0 140.7 2.8 ;
    END
  END s_vinj<1>
  PIN s_vinj<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 153.3 0.0 154.7 2.8 ;
    END
  END s_vinj<2>
  PIN s_gnd<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 167.3 0.0 168.7 2.8 ;
    END
  END s_gnd<0>
  PIN s_gnd<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 181.3 0.0 182.7 2.8 ;
    END
  END s_gnd<1>
  PIN s_gnd<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 195.3 0.0 196.7 2.8 ;
    END
  END s_gnd<2>
  PIN s_avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 209.3 0.0 210.7 2.8 ;
    END
  END s_avdd
  PIN s_s0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 223.3 0.0 224.7 2.8 ;
    END
  END s_s0
  PIN s_s1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 237.3 0.0 238.7 2.8 ;
    END
  END s_s1
  PIN s_s2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 251.3 0.0 252.7 2.8 ;
    END
  END s_s2
  PIN s_s3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 265.3 0.0 266.7 2.8 ;
    END
  END s_s3
  PIN s_s4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 279.3 0.0 280.7 2.8 ;
    END
  END s_s4
  PIN s_s5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 293.3 0.0 294.7 2.8 ;
    END
  END s_s5
  PIN s_s6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 307.3 0.0 308.7 2.8 ;
    END
  END s_s6
  PIN s_s7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 321.3 0.0 322.7 2.8 ;
    END
  END s_s7
  PIN s_s8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 335.3 0.0 336.7 2.8 ;
    END
  END s_s8
  PIN s_s9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 349.3 0.0 350.7 2.8 ;
    END
  END s_s9
  PIN s_s10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 363.3 0.0 364.7 2.8 ;
    END
  END s_s10
  PIN s_s11
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 377.3 0.0 378.7 2.8 ;
    END
  END s_s11
  PIN s_prog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 391.3 0.0 392.7 2.8 ;
    END
  END s_prog
  PIN s_run
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 405.3 0.0 406.7 2.8 ;
    END
  END s_run
  PIN s_vgsel
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 419.3 0.0 420.7 2.8 ;
    END
  END s_vgsel
  PIN w_cns0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 551.99 2.8 553.39 ;
    END
  END w_cns0
  PIN w_cns1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 537.99 2.8 539.39 ;
    END
  END w_cns1
  PIN w_cns2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 523.99 2.8 525.39 ;
    END
  END w_cns2
  PIN w_cns3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 509.99 2.8 511.39 ;
    END
  END w_cns3
  PIN w_vgrun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 495.99 2.8 497.39 ;
    END
  END w_vgrun
  PIN w_vtun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 481.99 2.8 483.39 ;
    END
  END w_vtun
  PIN w_vinj
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 467.99 2.8 469.39 ;
    END
  END w_vinj
  PIN w_gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 453.99 2.8 455.39 ;
    END
  END w_gnd
  PIN w_avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 439.99 2.8 441.39 ;
    END
  END w_avdd
  PIN w_drainbit3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 425.99 2.8 427.39 ;
    END
  END w_drainbit3
  PIN w_drainbit2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 411.99 2.8 413.39 ;
    END
  END w_drainbit2
  PIN w_drainbit1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 397.99 2.8 399.39 ;
    END
  END w_drainbit1
  PIN w_drainbit0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 383.99 2.8 385.39 ;
    END
  END w_drainbit0
  PIN w_s0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 369.99 2.8 371.39 ;
    END
  END w_s0
  PIN w_s1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 355.99 2.8 357.39 ;
    END
  END w_s1
  PIN w_s2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 341.99 2.8 343.39 ;
    END
  END w_s2
  PIN w_s3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 327.99 2.8 329.39 ;
    END
  END w_s3
  PIN w_s4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 313.99 2.8 315.39 ;
    END
  END w_s4
  PIN w_s5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 299.99 2.8 301.39 ;
    END
  END w_s5
  PIN w_s6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 285.99 2.8 287.39 ;
    END
  END w_s6
  PIN w_s7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 271.99 2.8 273.39 ;
    END
  END w_s7
  PIN w_s8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 257.99 2.8 259.39 ;
    END
  END w_s8
  PIN w_s9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 243.99 2.8 245.39 ;
    END
  END w_s9
  PIN w_s10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 229.99 2.8 231.39 ;
    END
  END w_s10
  PIN w_s11
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 215.99 2.8 217.39 ;
    END
  END w_s11
  PIN w_drainbit9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 201.99 2.8 203.39 ;
    END
  END w_drainbit9
  PIN w_drainbit8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 187.99 2.8 189.39 ;
    END
  END w_drainbit8
  PIN w_drainbit7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 173.99 2.8 175.39 ;
    END
  END w_drainbit7
  PIN w_drainbit6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 159.99 2.8 161.39 ;
    END
  END w_drainbit6
  PIN w_drainbit5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 145.99 2.8 147.39 ;
    END
  END w_drainbit5
  PIN w_drainbit4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 131.99 2.8 133.39 ;
    END
  END w_drainbit4
  PIN w_drainEN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 117.99 2.8 119.39 ;
    END
  END w_drainEN
END cab1

MACRO cab2
  PIN n_gateEN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 13.3 629.09 14.7 631.89 ;
    END
  END n_gateEN
  PIN n_programdrain
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 27.3 629.09 28.7 631.89 ;
    END
  END n_programdrain
  PIN n_rundrain
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 41.3 629.09 42.7 631.89 ;
    END
  END n_rundrain
  PIN n_cew0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 55.3 629.09 56.7 631.89 ;
    END
  END n_cew0
  PIN n_cew1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 69.3 629.09 70.7 631.89 ;
    END
  END n_cew1
  PIN n_cew2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 83.3 629.09 84.7 631.89 ;
    END
  END n_cew2
  PIN n_cew3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.3 629.09 98.7 631.89 ;
    END
  END n_cew3
  PIN n_vtun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 111.3 629.09 112.7 631.89 ;
    END
  END n_vtun
  PIN n_vinj<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 125.3 629.09 126.7 631.89 ;
    END
  END n_vinj<0>
  PIN n_vinj<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 139.3 629.09 140.7 631.89 ;
    END
  END n_vinj<1>
  PIN n_vinj<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 153.3 629.09 154.7 631.89 ;
    END
  END n_vinj<2>
  PIN n_gnd<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 167.3 629.09 168.7 631.89 ;
    END
  END n_gnd<0>
  PIN n_gnd<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 181.3 629.09 182.7 631.89 ;
    END
  END n_gnd<1>
  PIN n_gnd<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 195.3 629.09 196.7 631.89 ;
    END
  END n_gnd<2>
  PIN n_avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 209.3 629.09 210.7 631.89 ;
    END
  END n_avdd
  PIN n_s0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 223.3 629.09 224.7 631.89 ;
    END
  END n_s0
  PIN n_s1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 237.3 629.09 238.7 631.89 ;
    END
  END n_s1
  PIN n_s2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 251.3 629.09 252.7 631.89 ;
    END
  END n_s2
  PIN n_s3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 265.3 629.09 266.7 631.89 ;
    END
  END n_s3
  PIN n_s4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 279.3 629.09 280.7 631.89 ;
    END
  END n_s4
  PIN n_s5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 293.3 629.09 294.7 631.89 ;
    END
  END n_s5
  PIN n_s6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 307.3 629.09 308.7 631.89 ;
    END
  END n_s6
  PIN n_s7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 321.3 629.09 322.7 631.89 ;
    END
  END n_s7
  PIN n_s8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 335.3 629.09 336.7 631.89 ;
    END
  END n_s8
  PIN n_s9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 349.3 629.09 350.7 631.89 ;
    END
  END n_s9
  PIN n_s10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 363.3 629.09 364.7 631.89 ;
    END
  END n_s10
  PIN n_s11
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 377.3 629.09 378.7 631.89 ;
    END
  END n_s11
  PIN n_s12
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 391.3 629.09 392.7 631.89 ;
    END
  END n_s12
  PIN n_s13
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 405.3 629.09 406.7 631.89 ;
    END
  END n_s13
  PIN n_s14
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 419.3 629.09 420.7 631.89 ;
    END
  END n_s14
  PIN n_s15
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 433.3 629.09 434.7 631.89 ;
    END
  END n_s15
  PIN n_s16
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 447.3 629.09 448.7 631.89 ;
    END
  END n_s16
  PIN n_s17
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 461.3 629.09 462.7 631.89 ;
    END
  END n_s17
  PIN n_s18
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 475.3 629.09 476.7 631.89 ;
    END
  END n_s18
  PIN n_s19
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 489.3 629.09 490.7 631.89 ;
    END
  END n_s19
  PIN n_s20
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 503.3 629.09 504.7 631.89 ;
    END
  END n_s20
  PIN n_s21
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 517.3 629.09 518.7 631.89 ;
    END
  END n_s21
  PIN n_s22
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 531.3 629.09 532.7 631.89 ;
    END
  END n_s22
  PIN n_s23
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 545.3 629.09 546.7 631.89 ;
    END
  END n_s23
  PIN n_prog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 559.3 629.09 560.7 631.89 ;
    END
  END n_prog
  PIN n_run
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 573.3 629.09 574.7 631.89 ;
    END
  END n_run
  PIN n_vgsel
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 587.3 629.09 588.7 631.89 ;
    END
  END n_vgsel
  PIN e_cns0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 616.49 875.45 617.89 ;
    END
  END e_cns0
  PIN e_cns1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 602.49 875.45 603.89 ;
    END
  END e_cns1
  PIN e_cns2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 588.49 875.45 589.89 ;
    END
  END e_cns2
  PIN e_cns3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 574.49 875.45 575.89 ;
    END
  END e_cns3
  PIN e_vgrun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 560.49 875.45 561.89 ;
    END
  END e_vgrun
  PIN e_vtun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 546.49 875.45 547.89 ;
    END
  END e_vtun
  PIN e_vinj
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 532.49 875.45 533.89 ;
    END
  END e_vinj
  PIN e_gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 518.49 875.45 519.89 ;
    END
  END e_gnd
  PIN e_avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 504.49 875.45 505.89 ;
    END
  END e_avdd
  PIN e_drainbit4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 490.49 875.45 491.89 ;
    END
  END e_drainbit4
  PIN e_drainbit3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 476.49 875.45 477.89 ;
    END
  END e_drainbit3
  PIN e_drainbit2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 462.49 875.45 463.89 ;
    END
  END e_drainbit2
  PIN e_drainbit1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 448.49 875.45 449.89 ;
    END
  END e_drainbit1
  PIN e_drainbit0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 434.49 875.45 435.89 ;
    END
  END e_drainbit0
  PIN e_s0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 420.49 875.45 421.89 ;
    END
  END e_s0
  PIN e_s1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 406.49 875.45 407.89 ;
    END
  END e_s1
  PIN e_s2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 392.49 875.45 393.89 ;
    END
  END e_s2
  PIN e_s3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 378.49 875.45 379.89 ;
    END
  END e_s3
  PIN e_s4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 364.49 875.45 365.89 ;
    END
  END e_s4
  PIN e_s5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 350.49 875.45 351.89 ;
    END
  END e_s5
  PIN e_s6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 336.49 875.45 337.89 ;
    END
  END e_s6
  PIN e_s7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 322.49 875.45 323.89 ;
    END
  END e_s7
  PIN e_s8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 308.49 875.45 309.89 ;
    END
  END e_s8
  PIN e_s9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 294.49 875.45 295.89 ;
    END
  END e_s9
  PIN e_s10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 280.49 875.45 281.89 ;
    END
  END e_s10
  PIN e_s11
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 266.49 875.45 267.89 ;
    END
  END e_s11
  PIN e_s12
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 252.49 875.45 253.89 ;
    END
  END e_s12
  PIN e_s13
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 238.49 875.45 239.89 ;
    END
  END e_s13
  PIN e_s14
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 224.49 875.45 225.89 ;
    END
  END e_s14
  PIN e_s15
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 210.49 875.45 211.89 ;
    END
  END e_s15
  PIN e_s16
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 196.49 875.45 197.89 ;
    END
  END e_s16
  PIN e_s17
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 182.49 875.45 183.89 ;
    END
  END e_s17
  PIN e_s18
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 168.49 875.45 169.89 ;
    END
  END e_s18
  PIN e_s19
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 154.49 875.45 155.89 ;
    END
  END e_s19
  PIN e_s20
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 140.49 875.45 141.89 ;
    END
  END e_s20
  PIN e_s21
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 126.49 875.45 127.89 ;
    END
  END e_s21
  PIN e_s22
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 112.49 875.45 113.89 ;
    END
  END e_s22
  PIN e_s23
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 98.49 875.45 99.89 ;
    END
  END e_s23
  PIN e_drainbit10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 84.49 875.45 85.89 ;
    END
  END e_drainbit10
  PIN e_drainbit9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 70.49 875.45 71.89 ;
    END
  END e_drainbit9
  PIN e_drainbit8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 56.49 875.45 57.89 ;
    END
  END e_drainbit8
  PIN e_drainbit7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 42.49 875.45 43.89 ;
    END
  END e_drainbit7
  PIN e_drainbit6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 28.49 875.45 29.89 ;
    END
  END e_drainbit6
  PIN e_drainbit5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 14.49 875.45 15.89 ;
    END
  END e_drainbit5
  PIN e_drainEN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 872.65 0.49 875.45 1.89 ;
    END
  END e_drainEN
  PIN s_gateEN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 13.3 0.0 14.7 2.8 ;
    END
  END s_gateEN
  PIN s_programdrain
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 27.3 0.0 28.7 2.8 ;
    END
  END s_programdrain
  PIN s_rundrain
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 41.3 0.0 42.7 2.8 ;
    END
  END s_rundrain
  PIN s_cew0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 55.3 0.0 56.7 2.8 ;
    END
  END s_cew0
  PIN s_cew1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 69.3 0.0 70.7 2.8 ;
    END
  END s_cew1
  PIN s_cew2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 83.3 0.0 84.7 2.8 ;
    END
  END s_cew2
  PIN s_cew3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.3 0.0 98.7 2.8 ;
    END
  END s_cew3
  PIN s_vtun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 111.3 0.0 112.7 2.8 ;
    END
  END s_vtun
  PIN s_vinj<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 125.3 0.0 126.7 2.8 ;
    END
  END s_vinj<0>
  PIN s_vinj<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 139.3 0.0 140.7 2.8 ;
    END
  END s_vinj<1>
  PIN s_vinj<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 153.3 0.0 154.7 2.8 ;
    END
  END s_vinj<2>
  PIN s_gnd<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 167.3 0.0 168.7 2.8 ;
    END
  END s_gnd<0>
  PIN s_gnd<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 181.3 0.0 182.7 2.8 ;
    END
  END s_gnd<1>
  PIN s_gnd<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 195.3 0.0 196.7 2.8 ;
    END
  END s_gnd<2>
  PIN s_avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 209.3 0.0 210.7 2.8 ;
    END
  END s_avdd
  PIN s_s0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 223.3 0.0 224.7 2.8 ;
    END
  END s_s0
  PIN s_s1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 237.3 0.0 238.7 2.8 ;
    END
  END s_s1
  PIN s_s2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 251.3 0.0 252.7 2.8 ;
    END
  END s_s2
  PIN s_s3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 265.3 0.0 266.7 2.8 ;
    END
  END s_s3
  PIN s_s4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 279.3 0.0 280.7 2.8 ;
    END
  END s_s4
  PIN s_s5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 293.3 0.0 294.7 2.8 ;
    END
  END s_s5
  PIN s_s6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 307.3 0.0 308.7 2.8 ;
    END
  END s_s6
  PIN s_s7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 321.3 0.0 322.7 2.8 ;
    END
  END s_s7
  PIN s_s8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 335.3 0.0 336.7 2.8 ;
    END
  END s_s8
  PIN s_s9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 349.3 0.0 350.7 2.8 ;
    END
  END s_s9
  PIN s_s10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 363.3 0.0 364.7 2.8 ;
    END
  END s_s10
  PIN s_s11
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 377.3 0.0 378.7 2.8 ;
    END
  END s_s11
  PIN s_s12
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 391.3 0.0 392.7 2.8 ;
    END
  END s_s12
  PIN s_s13
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 405.3 0.0 406.7 2.8 ;
    END
  END s_s13
  PIN s_s14
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 419.3 0.0 420.7 2.8 ;
    END
  END s_s14
  PIN s_s15
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 433.3 0.0 434.7 2.8 ;
    END
  END s_s15
  PIN s_s16
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 447.3 0.0 448.7 2.8 ;
    END
  END s_s16
  PIN s_s17
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 461.3 0.0 462.7 2.8 ;
    END
  END s_s17
  PIN s_s18
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 475.3 0.0 476.7 2.8 ;
    END
  END s_s18
  PIN s_s19
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 489.3 0.0 490.7 2.8 ;
    END
  END s_s19
  PIN s_s20
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 503.3 0.0 504.7 2.8 ;
    END
  END s_s20
  PIN s_s21
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 517.3 0.0 518.7 2.8 ;
    END
  END s_s21
  PIN s_s22
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 531.3 0.0 532.7 2.8 ;
    END
  END s_s22
  PIN s_s23
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 545.3 0.0 546.7 2.8 ;
    END
  END s_s23
  PIN s_prog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 559.3 0.0 560.7 2.8 ;
    END
  END s_prog
  PIN s_run
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 573.3 0.0 574.7 2.8 ;
    END
  END s_run
  PIN s_vgsel
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 587.3 0.0 588.7 2.8 ;
    END
  END s_vgsel
  PIN w_cns0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 616.49 2.8 617.89 ;
    END
  END w_cns0
  PIN w_cns1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 602.49 2.8 603.89 ;
    END
  END w_cns1
  PIN w_cns2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 588.49 2.8 589.89 ;
    END
  END w_cns2
  PIN w_cns3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 574.49 2.8 575.89 ;
    END
  END w_cns3
  PIN w_vgrun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 560.49 2.8 561.89 ;
    END
  END w_vgrun
  PIN w_vtun
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 546.49 2.8 547.89 ;
    END
  END w_vtun
  PIN w_vinj
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 532.49 2.8 533.89 ;
    END
  END w_vinj
  PIN w_gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 518.49 2.8 519.89 ;
    END
  END w_gnd
  PIN w_avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 504.49 2.8 505.89 ;
    END
  END w_avdd
  PIN w_drainbit4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 490.49 2.8 491.89 ;
    END
  END w_drainbit4
  PIN w_drainbit3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 476.49 2.8 477.89 ;
    END
  END w_drainbit3
  PIN w_drainbit2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 462.49 2.8 463.89 ;
    END
  END w_drainbit2
  PIN w_drainbit1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 448.49 2.8 449.89 ;
    END
  END w_drainbit1
  PIN w_drainbit0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 434.49 2.8 435.89 ;
    END
  END w_drainbit0
  PIN w_s0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 420.49 2.8 421.89 ;
    END
  END w_s0
  PIN w_s1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 406.49 2.8 407.89 ;
    END
  END w_s1
  PIN w_s2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 392.49 2.8 393.89 ;
    END
  END w_s2
  PIN w_s3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 378.49 2.8 379.89 ;
    END
  END w_s3
  PIN w_s4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 364.49 2.8 365.89 ;
    END
  END w_s4
  PIN w_s5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 350.49 2.8 351.89 ;
    END
  END w_s5
  PIN w_s6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 336.49 2.8 337.89 ;
    END
  END w_s6
  PIN w_s7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 322.49 2.8 323.89 ;
    END
  END w_s7
  PIN w_s8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 308.49 2.8 309.89 ;
    END
  END w_s8
  PIN w_s9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 294.49 2.8 295.89 ;
    END
  END w_s9
  PIN w_s10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 280.49 2.8 281.89 ;
    END
  END w_s10
  PIN w_s11
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 266.49 2.8 267.89 ;
    END
  END w_s11
  PIN w_s12
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 252.49 2.8 253.89 ;
    END
  END w_s12
  PIN w_s13
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 238.49 2.8 239.89 ;
    END
  END w_s13
  PIN w_s14
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 224.49 2.8 225.89 ;
    END
  END w_s14
  PIN w_s15
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 210.49 2.8 211.89 ;
    END
  END w_s15
  PIN w_s16
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 196.49 2.8 197.89 ;
    END
  END w_s16
  PIN w_s17
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 182.49 2.8 183.89 ;
    END
  END w_s17
  PIN w_s18
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 168.49 2.8 169.89 ;
    END
  END w_s18
  PIN w_s19
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 154.49 2.8 155.89 ;
    END
  END w_s19
  PIN w_s20
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 140.49 2.8 141.89 ;
    END
  END w_s20
  PIN w_s21
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 126.49 2.8 127.89 ;
    END
  END w_s21
  PIN w_s22
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 112.49 2.8 113.89 ;
    END
  END w_s22
  PIN w_s23
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 98.49 2.8 99.89 ;
    END
  END w_s23
  PIN w_drainbit10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 84.49 2.8 85.89 ;
    END
  END w_drainbit10
  PIN w_drainbit9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 70.49 2.8 71.89 ;
    END
  END w_drainbit9
  PIN w_drainbit8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 56.49 2.8 57.89 ;
    END
  END w_drainbit8
  PIN w_drainbit7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 42.49 2.8 43.89 ;
    END
  END w_drainbit7
  PIN w_drainbit6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 28.49 2.8 29.89 ;
    END
  END w_drainbit6
  PIN w_drainbit5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 14.49 2.8 15.89 ;
    END
  END w_drainbit5
  PIN w_drainEN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 0.49 2.8 1.89 ;
    END
  END w_drainEN
END cab2

END LIBRARY