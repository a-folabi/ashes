module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(7), .GND_b_1_row_4(net2030[0:7]), .Vs_b_0_row_4(net124[0:7]), .Vs_b_1_row_4(net125[0:7]), .VINJ_b_1_row_4(net2037[0:7]), .Vsel_b_0_row_4(net1995[0:7]), .Vsel_b_1_row_4(net1996[0:7]), .Vg_b_0_row_4(net2009[0:7]), .Vg_b_1_row_4(net2010[0:7]), .VTUN_brow_4(net2023[0:7]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(17), .matrix_row(5), .matrix_col(9), .GND_b_1_row_4(net2073[0:9]), .Vs_b_0_row_4(net285[0:9]), .Vs_b_1_row_4(net286[0:9]), .VINJ_b_1_row_4(net2072[0:9]), .Vsel_b_0_row_4(net2074[0:9]), .Vsel_b_1_row_4(net2076[0:9]), .Vg_b_0_row_4(net304[0:9]), .Vg_b_1_row_4(net305[0:9]), .VTUN_brow_4(net2071[0:9]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(26), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2050[0:1]), .Vsel_b_0_row_4(net2053[0:1]), .Vsel_b_1_row_4(net2054[0:1]), .Vg_b_0_row_4(net2055[0:1]), .Vg_b_1_row_4(net2056[0:1]), .VTUN_brow_4(net2051[0:1]), .GND_b_1_row_4(net2052[0:1]));
	S_BLOCK_BUFFER I__4 (.island_num(0), .row(0), .col(8), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__5 (.island_num(0), .row(0), .col(9), .matrix_row(4), .matrix_col(1));
	S_BLOCK_CONN_PINS I__6 (.island_num(0), .row(4), .col(9), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__7 (.island_num(0), .row(0), .col(10), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__8 (.island_num(0), .row(3), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__9 (.island_num(0), .row(4), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__10 (.island_num(0), .row(0), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_CONN_PINS I__11 (.island_num(0), .row(2), .col(11), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__12 (.island_num(0), .row(3), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__13 (.island_num(0), .row(0), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_CONN_PINS I__14 (.island_num(0), .row(1), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__15 (.island_num(0), .row(2), .col(12), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__16 (.island_num(0), .row(0), .col(13), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__17 (.island_num(0), .row(1), .col(13), .matrix_row(4), .matrix_col(1));
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2057[0:1]), .Vsel_b_0_row_4(net2060[0:1]), .Vsel_b_1_row_4(net2061[0:1]), .Vg_b_0_row_4(net2062[0:1]), .Vg_b_1_row_4(net2063[0:1]), .VTUN_brow_4(net2058[0:1]), .GND_b_1_row_4(net2059[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2064[0:1]), .Vsel_b_0_row_4(net2067[0:1]), .Vsel_b_1_row_4(net2068[0:1]), .Vg_b_0_row_4(net2069[0:1]), .Vg_b_1_row_4(net2070[0:1]), .VTUN_brow_4(net2065[0:1]), .GND_b_1_row_4(net2066[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(6), .decode_n0_RUN_OUT_0_(net2144), .decode_n0_RUN_OUT_1_(net2145), .decode_n0_RUN_OUT_2_(net2150), .decode_n0_RUN_OUT_3_(net2151), .decode_n1_RUN_OUT_0_(net2156), .decode_n1_RUN_OUT_1_(net2157), .decode_n1_RUN_OUT_2_(net2162), .decode_n1_RUN_OUT_3_(net2163), .decode_n2_RUN_OUT_0_(net2168), .decode_n2_RUN_OUT_1_(net2169), .decode_n2_RUN_OUT_2_(net2174), .decode_n2_RUN_OUT_3_(net2175), .decode_n3_RUN_OUT_0_(net2180), .decode_n3_RUN_OUT_1_(net2181), .decode_n3_RUN_OUT_2_(net2186), .decode_n3_RUN_OUT_3_(net2187), .decode_n4_RUN_OUT_2_(net2192), .decode_n4_RUN_OUT_3_(net2193), .decode_n5_RUN_OUT_0_(net2198), .decode_n5_RUN_OUT_1_(net2199), .decode_n5_RUN_OUT_2_(net2204), .decode_n5_RUN_OUT_3_(net2205), .decode_n6_RUN_OUT_0_(net2210), .decode_n6_RUN_OUT_1_(net2211), .decode_n6_RUN_OUT_2_(net2216), .decode_n6_RUN_OUT_3_(net2217), .decode_n7_RUN_OUT_0_(net2222), .decode_n7_RUN_OUT_1_(net2223), .decode_n7_RUN_OUT_2_(net2228), .decode_n7_RUN_OUT_3_(net2229), .decode_n8_RUN_OUT_0_(net2234), .decode_n8_RUN_OUT_1_(net2235), .decode_n8_RUN_OUT_2_(net2240), .decode_n8_RUN_OUT_3_(net2241), .decode_n9_RUN_OUT_0_(net2246), .decode_n9_RUN_OUT_1_(net2247), .decode_n9_RUN_OUT_2_(net2252), .decode_n9_RUN_OUT_3_(net2253), .decode_n0_OUT_0_(net2142), .decode_n0_OUT_1_(net2143), .decode_n0_OUT_2_(net2148), .decode_n0_OUT_3_(net2149), .decode_n1_OUT_0_(net2154), .decode_n1_OUT_1_(net2155), .decode_n1_OUT_2_(net2160), .decode_n1_OUT_3_(net2161), .decode_n2_OUT_0_(net2166), .decode_n2_OUT_1_(net2167), .decode_n2_OUT_2_(net2172), .decode_n2_OUT_3_(net2173), .decode_n3_OUT_0_(net2178), .decode_n3_OUT_1_(net2179), .decode_n3_OUT_2_(net2184), .decode_n3_OUT_3_(net2185), .decode_n4_OUT_2_(net2190), .decode_n4_OUT_3_(net2191), .decode_n5_OUT_0_(net2196), .decode_n5_OUT_1_(net2197), .decode_n5_OUT_2_(net2202), .decode_n5_OUT_3_(net2203), .decode_n6_OUT_0_(net2208), .decode_n6_OUT_1_(net2209), .decode_n6_OUT_2_(net2214), .decode_n6_OUT_3_(net2215), .decode_n7_OUT_0_(net2220), .decode_n7_OUT_1_(net2221), .decode_n7_OUT_2_(net2226), .decode_n7_OUT_3_(net2227), .decode_n8_OUT_0_(net2232), .decode_n8_OUT_1_(net2233), .decode_n8_OUT_2_(net2238), .decode_n8_OUT_3_(net2239), .decode_n9_OUT_0_(net2244), .decode_n9_OUT_1_(net2245), .decode_n9_OUT_2_(net2250), .decode_n9_OUT_3_(net2251), .decode_n0_VINJ_b_0_(net2140), .decode_n0_VINJ_b_1_(net2146), .decode_n1_VINJ_b_0_(net2152), .decode_n1_VINJ_b_1_(net2158), .decode_n2_VINJ_b_0_(net2164), .decode_n2_VINJ_b_1_(net2170), .decode_n3_VINJ_b_0_(net2176), .decode_n3_VINJ_b_1_(net2182), .decode_n4_VINJ_b_1_(net2188), .decode_n5_VINJ_b_0_(net2194), .decode_n5_VINJ_b_1_(net2200), .decode_n6_VINJ_b_0_(net2206), .decode_n6_VINJ_b_1_(net2212), .decode_n7_VINJ_b_0_(net2218), .decode_n7_VINJ_b_1_(net2224), .decode_n8_VINJ_b_0_(net2230), .decode_n8_VINJ_b_1_(net2236), .decode_n9_VINJ_b_0_(net2242), .decode_n9_VINJ_b_1_(net2248), .decode_n0_GND_b_0_(net2141), .decode_n0_GND_b_1_(net2147), .decode_n1_GND_b_0_(net2153), .decode_n1_GND_b_1_(net2159), .decode_n2_GND_b_0_(net2165), .decode_n2_GND_b_1_(net2171), .decode_n3_GND_b_0_(net2177), .decode_n3_GND_b_1_(net2183), .decode_n4_GND_b_1_(net2189), .decode_n5_GND_b_0_(net2195), .decode_n5_GND_b_1_(net2201), .decode_n6_GND_b_0_(net2207), .decode_n6_GND_b_1_(net2213), .decode_n7_GND_b_0_(net2219), .decode_n7_GND_b_1_(net2225), .decode_n8_GND_b_0_(net2231), .decode_n8_GND_b_1_(net2237), .decode_n9_GND_b_0_(net2243), .decode_n9_GND_b_1_(net2249));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(26), .switch_n0_VPWR_0_(net2144), .switch_n0_VPWR_1_(net2145), .switch_n1_VPWR_0_(net2150), .switch_n1_VPWR_1_(net2151), .switch_n2_VPWR_0_(net2156), .switch_n2_VPWR_1_(net2157), .switch_n3_VPWR_0_(net2162), .switch_n3_VPWR_1_(net2163), .switch_n4_VPWR_0_(net2168), .switch_n4_VPWR_1_(net2169), .switch_n5_VPWR_0_(net2174), .switch_n5_VPWR_1_(net2175), .switch_n6_VPWR_0_(net2180), .switch_n6_VPWR_1_(net2181), .switch_n7_VPWR_0_(net2186), .switch_n7_VPWR_1_(net2187), .switch_n14_VPWR_0_(net2192), .switch_n14_VPWR_1_(net2193), .switch_n16_VPWR_0_(net2198), .switch_n16_VPWR_1_(net2199), .switch_n17_VPWR_0_(net2204), .switch_n17_VPWR_1_(net2205), .switch_n18_VPWR_0_(net2210), .switch_n18_VPWR_1_(net2211), .switch_n19_VPWR_0_(net2216), .switch_n19_VPWR_1_(net2217), .switch_n20_VPWR_0_(net2222), .switch_n20_VPWR_1_(net2223), .switch_n21_VPWR_0_(net2228), .switch_n21_VPWR_1_(net2229), .switch_n22_VPWR_0_(net2234), .switch_n22_VPWR_1_(net2235), .switch_n23_VPWR_0_(net2240), .switch_n23_VPWR_1_(net2241), .switch_n24_VPWR_0_(net2246), .switch_n24_VPWR_1_(net2247), .switch_n25_VPWR_0_(net2252), .switch_n25_VPWR_1_(net2253), .switch_n0_GND_T(net2141), .switch_n1_GND_T(net2147), .switch_n2_GND_T(net2153), .switch_n3_GND_T(net2159), .switch_n4_GND_T(net2165), .switch_n5_GND_T(net2171), .switch_n6_GND_T(net2177), .switch_n7_GND_T(net2183), .switch_n14_GND_T(net2189), .switch_n16_GND_T(net2195), .switch_n17_GND_T(net2201), .switch_n18_GND_T(net2207), .switch_n19_GND_T(net2213), .switch_n20_GND_T(net2219), .switch_n21_GND_T(net2225), .switch_n22_GND_T(net2231), .switch_n23_GND_T(net2237), .switch_n24_GND_T(net2243), .switch_n25_GND_T(net2249), .switch_n0_decode_0_(net2142), .switch_n0_decode_1_(net2143), .switch_n1_decode_0_(net2148), .switch_n1_decode_1_(net2149), .switch_n2_decode_0_(net2154), .switch_n2_decode_1_(net2155), .switch_n3_decode_0_(net2160), .switch_n3_decode_1_(net2161), .switch_n4_decode_0_(net2166), .switch_n4_decode_1_(net2167), .switch_n5_decode_0_(net2172), .switch_n5_decode_1_(net2173), .switch_n6_decode_0_(net2178), .switch_n6_decode_1_(net2179), .switch_n7_decode_0_(net2184), .switch_n7_decode_1_(net2185), .switch_n14_decode_0_(net2190), .switch_n14_decode_1_(net2191), .switch_n16_decode_0_(net2196), .switch_n16_decode_1_(net2197), .switch_n17_decode_0_(net2202), .switch_n17_decode_1_(net2203), .switch_n18_decode_0_(net2208), .switch_n18_decode_1_(net2209), .switch_n19_decode_0_(net2214), .switch_n19_decode_1_(net2215), .switch_n20_decode_0_(net2220), .switch_n20_decode_1_(net2221), .switch_n21_decode_0_(net2226), .switch_n21_decode_1_(net2227), .switch_n22_decode_0_(net2232), .switch_n22_decode_1_(net2233), .switch_n23_decode_0_(net2238), .switch_n23_decode_1_(net2239), .switch_n24_decode_0_(net2244), .switch_n24_decode_1_(net2245), .switch_n25_decode_0_(net2250), .switch_n25_decode_1_(net2251), .switch_n0_VINJ_T(net2140), .switch_n1_VINJ_T(net2146), .switch_n2_VINJ_T(net2152), .switch_n3_VINJ_T(net2158), .switch_n4_VINJ_T(net2164), .switch_n5_VINJ_T(net2170), .switch_n6_VINJ_T(net2176), .switch_n7_VINJ_T(net2182), .switch_n14_VINJ_T(net2188), .switch_n16_VINJ_T(net2194), .switch_n17_VINJ_T(net2200), .switch_n18_VINJ_T(net2206), .switch_n19_VINJ_T(net2212), .switch_n20_VINJ_T(net2218), .switch_n21_VINJ_T(net2224), .switch_n22_VINJ_T(net2230), .switch_n23_VINJ_T(net2236), .switch_n24_VINJ_T(net2242), .switch_n25_VINJ_T(net2248));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch));
	none switch_ind(.island_num(0), .direction(horizontal), .col(8));
	none switch_ind(.island_num(0), .direction(horizontal), .col(9));
	none switch_ind(.island_num(0), .direction(horizontal), .col(10));
	none switch_ind(.island_num(0), .direction(horizontal), .col(11));
	none switch_ind(.island_num(0), .direction(horizontal), .col(12));
	none switch_ind(.island_num(0), .direction(horizontal), .col(13));
	none switch_ind(.island_num(0), .direction(horizontal), .col(15));


	/* Island 1 */
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__0 (.island_num(1), .row(0), .col(0), .matrix_row(1), .matrix_col(8));
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(7), .matrix_col(8), .GND_b_0_row_6(net1138[0:8]), .GND_b_1_row_6(net1139[0:8]), .Vs_b_0_row_6(net1148[0:8]), .Vs_b_1_row_6(net1149[0:8]), .VINJ_b_0_row_6(net1152[0:8]), .VINJ_b_1_row_6(net1153[0:8]), .Vsel_b_0_row_6(net1156[0:8]), .Vsel_b_1_row_6(net1157[0:8]), .Vg_b_0_row_6(net1160[0:8]), .Vg_b_1_row_6(net1161[0:8]), .VTUN_brow_6(net1164[0:8]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(8), .matrix_row(6), .matrix_col(10));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(7), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1895), .P_1_row_0(net1896), .A_0_row_0(net1897), .A_1_row_0(net1898), .A_2_row_0(net1899), .A_3_row_0(net1900));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1908), .P_1_row_0(net1909), .A_0_row_0(net1910), .A_1_row_0(net1911), .A_2_row_0(net1912), .A_3_row_0(net1913));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1926), .P_1_row_0(net1927), .A_0_row_0(net1928), .A_1_row_0(net1929), .A_2_row_0(net1930), .A_3_row_0(net1931));
	TSMC350nm_4TGate_ST_BMatrix_NoSwitch I__8 (.island_num(1), .row(3), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1944), .P_1_row_0(net1945), .P_2_row_0(net1946), .P_3_row_0(net1947), .A_0_row_0(net1948), .A_1_row_0(net1949), .A_2_row_0(net1950), .A_3_row_0(net1951));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1963), .P_1_row_0(net1964), .P_2_row_0(net1965), .P_3_row_0(net1966), .A_0_row_0(net1967), .A_1_row_0(net1968));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1978), .A_1_row_0(net1979), .A_2_row_0(net1980), .A_3_row_0(net1981));
	TSMC350nm_4TGate_ST_BMatrix I__11 (.island_num(1), .row(6), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1985), .A_1_row_0(net1986), .A_2_row_0(net1987), .A_3_row_0(net1988));
	TSMC350nm_4TGate_ST_BMatrix I__12 (.island_num(1), .row(7), .col(18), .matrix_row(1), .matrix_col(1));
	TSMC350nm_OutMtrx_IndrctSwcs I__13 (.island_num(1), .row(9), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__14 (.island_num(1), .row(10), .col(8), .matrix_row(2), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__15 (.island_num(1), .row(10), .col(18), .matrix_row(2), .matrix_col(1));
	TSMC350nm_TA2Cell_Weak cab_device_16 (.island_num(1), .row(2), .col(19), .VD_P_0_(net1895), .VD_P_1_(net1896), .VIN1_PLUS(net1897), .VIN1_MINUS(net1898), .VIN2_PLUS(net1899), .VIN2_MINUS(net1900), .OUTPUT_0_(net1901[0]), .OUTPUT_1_(net1902[0]), .Vsel_0_(net1972), .Vsel_1_(net1973), .RUN(net1903), .Vg_0_(net1974), .Vg_1_(net1975), .PROG(net1904), .VTUN(net1905), .VINJ(net1906), .GND(net1907), .VPWR(net2317[0]), .Vsel_b_0_(net1916), .Vsel_b_1_(net1917), .RUN_b(net1918), .Vg_b_0_(net1919), .Vg_b_1_(net1920), .PROG_b(net1921), .VTUN_b(net1922), .VINJ_b(net1923), .GND_b(net1924), .VPWR_b(net1925));
	TSMC350nm_TA2Cell_Weak cab_device_17 (.island_num(1), .row(3), .col(19), .VD_P_0_(net1908), .VD_P_1_(net1909), .VIN1_PLUS(net1910), .VIN1_MINUS(net1911), .VIN2_PLUS(net1912), .VIN2_MINUS(net1913), .OUTPUT_0_(net1914[0]), .OUTPUT_1_(net1915[0]), .Vsel_0_(net1916), .Vsel_1_(net1917), .RUN(net1918), .Vg_0_(net1919), .Vg_1_(net1920), .PROG(net1921), .VTUN(net1922), .VINJ(net1923), .GND(net1924), .VPWR(net1925), .Vsel_b_0_(net1934), .Vsel_b_1_(net1935), .RUN_b(net1936), .Vg_b_0_(net1937), .Vg_b_1_(net1938), .PROG_b(net1939), .VTUN_b(net1940), .VINJ_b(net1941), .GND_b(net1942), .VPWR_b(net1943));
	TSMC350nm_TA2Cell_Strong cab_device_18 (.island_num(1), .row(4), .col(19), .VD_P_0_(net1926), .VD_P_1_(net1927), .VIN1_PLUS(net1928), .VIN1_MINUS(net1929), .VIN2_PLUS(net1930), .VIN2_MINUS(net1931), .OUTPUT_0_(net1932[0]), .OUTPUT_1_(net1933[0]), .Vsel_0_(net1934), .Vsel_1_(net1935), .RUN(net1936), .Vg_0_(net1937), .Vg_1_(net1938), .PROG(net1939), .VTUN(net1940), .VINJ(net1941), .GND(net1942), .VPWR(net1943), .Vg_b_0_(net1959), .PROG_b(net1962), .VTUN_b(net1960), .VINJ_b(net1958), .GND_b(net1961));
	TSMC350nm_4WTA_IndirectProg cab_device_19 (.island_num(1), .row(5), .col(19), .VD_P_0_(net1944), .VD_P_1_(net1945), .VD_P_2_(net1946), .VD_P_3_(net1947), .Iin_0_(net1948), .Iin_1_(net1949), .Iin_2_(net1950), .Iin_3_(net1951), .Vout_0_(net1952[0]), .Vout_1_(net1953[0]), .Vout_2_(net1954[0]), .Vout_3_(net1955[0]), .Vmid(net1956[0]), .Vbias(net1957[0]), .Vsel(net1972), .Vs(net2317[0]), .VINJ(net1958), .Vg(net1959), .VTUN(net1960), .GND(net1961), .PROG(net1962), .VINJ_b(net1971), .VTUN_b(net1977), .GND_b(net1976));
	TSMC350nm_Cap_Bank cab_device_20 (.island_num(1), .row(6), .col(19), .VD_P_0_(net1963), .VD_P_1_(net1964), .VD_P_2_(net1965), .VD_P_3_(net1966), .VIN_0_(net1967), .VIN_1_(net1968), .OUT_0_(net1969[0]), .OUT_1_(net1970[0]), .VINJ(net1971), .Vsel_0_(net1972), .Vsel_1_(net1973), .Vg_0_(net1974), .Vg_1_(net1975), .GND(net1976), .VTUN(net1977), .GND_b(net1984));
	TSMC350nm_NandPfets cab_device_21 (.island_num(1), .row(7), .col(19), .GATE_N(net1978), .SOURCE_N(net1979), .GATE_P(net1980), .SOURCE_P(net1981), .DRAIN_N(net1982[0]), .DRAIN_P(net1983[0]), .VPWR(net2317[0]), .GND(net1984), .VPWR_b(net1992), .GND_b(net1993));
	TSMC350nm_TGate_2nMirror cab_device_22 (.island_num(1), .row(8), .col(19), .IN_CM_0_(net1985), .IN_CM_1_(net1986), .SelN(net1987), .IN_TG(net1988), .OUT_CM_0_(net1989[0]), .OUT_CM_1_(net1990[0]), .OUT_TG(net1991[0]), .VPWR(net1992), .GND(net1993));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(1), .direction(vertical), .num(12), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(12), .type(prog_switch), .switch_n8_PR_3_(net2318[0]));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(20), .switch_n0_Input_0_(net1994), .switch_n0_Input_1_(net2030[0]), .switch_n1_Input_0_(net124[1]), .switch_n1_Input_1_(net125[1]), .switch_n2_Input_0_(net124[2]), .switch_n2_Input_1_(net125[2]), .switch_n3_Input_0_(net124[3]), .switch_n3_Input_1_(net125[3]), .switch_n4_Input_0_(net285[0]), .switch_n4_Input_1_(net286[0]), .switch_n5_Input_0_(net285[1]), .switch_n5_Input_1_(net286[1]), .switch_n6_Input_0_(net285[2]), .switch_n6_Input_1_(net286[2]), .switch_n7_Input_0_(net285[3]), .switch_n7_Input_1_(net286[3]), .switch_n8_Input_0_(net2316[0]), .switch_n8_Input_1_(net1901[0]), .switch_n9_Input_0_(net1902[0]), .switch_n9_Input_1_(net1914[0]), .switch_n10_Input_0_(net1915[0]), .switch_n10_Input_1_(net1932[0]), .switch_n11_Input_0_(net1933[0]), .switch_n11_Input_1_(net1952[0]), .switch_n12_Input_0_(net1953[0]), .switch_n12_Input_1_(net1954[0]), .switch_n13_Input_0_(net1955[0]), .switch_n13_Input_1_(net1956[0]), .switch_n14_Input_0_(net1957[0]), .switch_n14_Input_1_(net1969[0]), .switch_n15_Input_0_(net1970[0]), .switch_n15_Input_1_(net1982[0]), .switch_n16_Input_0_(net1983[0]), .switch_n16_Input_1_(net1989[0]), .switch_n17_Input_0_(net1990[0]), .switch_n17_Input_1_(net1991[0]), .switch_n0_GND(net2030[0]), .switch_n1_GND(net2030[1]), .switch_n2_GND(net2030[2]), .switch_n3_GND(net2030[3]), .switch_n4_GND(net2030[4]), .switch_n5_GND(net2030[5]), .switch_n6_GND(net2030[6]), .switch_n7_GND(net2052[0]), .switch_n8_GND(net2059[0]), .switch_n9_GND(net2066[0]), .switch_n10_GND(net2073[0]), .switch_n11_GND(net2073[1]), .switch_n12_GND(net2073[2]), .switch_n13_GND(net2073[3]), .switch_n14_GND(net2073[4]), .switch_n15_GND(net2073[5]), .switch_n16_GND(net2073[6]), .switch_n17_GND(net2073[7]), .switch_n0_Vsel_0_(net1995[0]), .switch_n0_Vsel_1_(net1996[0]), .switch_n1_Vsel_0_(net1995[1]), .switch_n1_Vsel_1_(net1996[1]), .switch_n2_Vsel_0_(net1995[2]), .switch_n2_Vsel_1_(net1996[2]), .switch_n3_Vsel_0_(net1995[3]), .switch_n3_Vsel_1_(net1996[3]), .switch_n4_Vsel_0_(net1995[4]), .switch_n4_Vsel_1_(net1996[4]), .switch_n5_Vsel_0_(net1995[5]), .switch_n5_Vsel_1_(net1996[5]), .switch_n6_Vsel_0_(net1995[6]), .switch_n6_Vsel_1_(net1996[6]), .switch_n7_Vsel_0_(net2054[0]), .switch_n7_Vsel_1_(net2053[0]), .switch_n8_Vsel_0_(net2061[0]), .switch_n8_Vsel_1_(net2060[0]), .switch_n9_Vsel_0_(net2068[0]), .switch_n9_Vsel_1_(net2067[0]), .switch_n10_Vsel_0_(net2074[0]), .switch_n10_Vsel_1_(net2076[0]), .switch_n11_Vsel_0_(net2074[1]), .switch_n11_Vsel_1_(net2076[1]), .switch_n12_Vsel_0_(net2074[2]), .switch_n12_Vsel_1_(net2076[2]), .switch_n13_Vsel_0_(net2074[3]), .switch_n13_Vsel_1_(net2076[3]), .switch_n14_Vsel_0_(net2074[4]), .switch_n14_Vsel_1_(net2076[4]), .switch_n15_Vsel_0_(net2074[5]), .switch_n15_Vsel_1_(net2076[5]), .switch_n16_Vsel_0_(net2074[6]), .switch_n16_Vsel_1_(net2076[6]), .switch_n17_Vsel_0_(net2074[7]), .switch_n17_Vsel_1_(net2076[7]), .switch_n0_Vg_global_0_(net2009[0]), .switch_n0_Vg_global_1_(net2010[0]), .switch_n1_Vg_global_0_(net2009[1]), .switch_n1_Vg_global_1_(net2010[1]), .switch_n2_Vg_global_0_(net2009[2]), .switch_n2_Vg_global_1_(net2010[2]), .switch_n3_Vg_global_0_(net2009[3]), .switch_n3_Vg_global_1_(net2010[3]), .switch_n4_Vg_global_0_(net2009[4]), .switch_n4_Vg_global_1_(net2010[4]), .switch_n5_Vg_global_0_(net2009[5]), .switch_n5_Vg_global_1_(net2010[5]), .switch_n6_Vg_global_0_(net2009[6]), .switch_n6_Vg_global_1_(net2010[6]), .switch_n7_Vg_global_0_(net2056[0]), .switch_n7_Vg_global_1_(net2055[0]), .switch_n8_Vg_global_0_(net2063[0]), .switch_n8_Vg_global_1_(net2062[0]), .switch_n9_Vg_global_0_(net2070[0]), .switch_n9_Vg_global_1_(net2069[0]), .switch_n10_Vg_global_0_(net304[0]), .switch_n10_Vg_global_1_(net305[0]), .switch_n11_Vg_global_0_(net304[1]), .switch_n11_Vg_global_1_(net305[1]), .switch_n12_Vg_global_0_(net304[2]), .switch_n12_Vg_global_1_(net305[2]), .switch_n13_Vg_global_0_(net304[3]), .switch_n13_Vg_global_1_(net305[3]), .switch_n14_Vg_global_0_(net304[4]), .switch_n14_Vg_global_1_(net305[4]), .switch_n15_Vg_global_0_(net304[5]), .switch_n15_Vg_global_1_(net305[5]), .switch_n16_Vg_global_0_(net304[6]), .switch_n16_Vg_global_1_(net305[6]), .switch_n17_Vg_global_0_(net304[7]), .switch_n17_Vg_global_1_(net305[7]), .switch_n0_VTUN(net2023[0]), .switch_n1_VTUN(net2023[1]), .switch_n2_VTUN(net2023[2]), .switch_n3_VTUN(net2023[3]), .switch_n4_VTUN(net2023[4]), .switch_n5_VTUN(net2023[5]), .switch_n6_VTUN(net2023[6]), .switch_n7_VTUN(net2051[0]), .switch_n8_VTUN(net2058[0]), .switch_n9_VTUN(net2065[0]), .switch_n10_VTUN(net2071[0]), .switch_n11_VTUN(net2071[1]), .switch_n12_VTUN(net2071[2]), .switch_n13_VTUN(net2071[3]), .switch_n14_VTUN(net2071[4]), .switch_n15_VTUN(net2071[5]), .switch_n16_VTUN(net2071[6]), .switch_n17_VTUN(net2071[7]), .switch_n0_VINJ(net2037[0]), .switch_n1_VINJ(net2037[1]), .switch_n2_VINJ(net2037[2]), .switch_n3_VINJ(net2037[3]), .switch_n4_VINJ(net2037[4]), .switch_n5_VINJ(net2037[5]), .switch_n6_VINJ(net2037[6]), .switch_n7_VINJ(net2050[0]), .switch_n8_VINJ(net2057[0]), .switch_n9_VINJ(net2064[0]), .switch_n10_VINJ(net2072[0]), .switch_n11_VINJ(net2072[1]), .switch_n12_VINJ(net2072[2]), .switch_n13_VINJ(net2072[3]), .switch_n14_VINJ(net2072[4]), .switch_n15_VINJ(net2072[5]), .switch_n16_VINJ(net2072[6]), .switch_n17_VINJ(net2072[7]));
	none switch_ind(.island_num(1), .direction(horizontal), .col(18));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(19), .VPWR_0_(net1994), .VPWR_1_(net1994), .GND_T(net2073[8]), .VTUN_T(net2071[8]), .decode_0_(net2074[8]), .decode_1_(net2076[8]), .VINJ_T(net2072[8]), .GND(net1907), .CTRL_B_0_(net1972), .CTRL_B_1_(net1973), .run_r(net1903), .prog_r(net1904), .Vg_0_(net1974), .Vg_1_(net1975), .VTUN(net1905), .VINJ(net1906), .VDD_1_(net2317[0]));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net1148[0:6]), .out_1_row_0(net1149[0:6]), .VINJ_0_row_0(net1152[0:6]), .VINJ_1_row_0(net1153[0:6]), .Vsel_0_row_0(net1156[0:6]), .Vsel_1_row_0(net1157[0:6]), .Vg_0_row_0(net1160[0:6]), .Vg_1_row_0(net1161[0:6]), .GNDrow_0(net1138[0:6]), .VTUNrow_0(net1164[0:6]), .Dcol_0(net124[6:7]), .CLKcol_0(net125[6:7]), .Qcol_5(net125[6:7]), .comcol_0(net2316[0:1]), .VDDcol_0(net2317[0:1]), .Vd_Pcol_0(net2318[0:1]));

 	/*Programming Mux */ 

 endmodule