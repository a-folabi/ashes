module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(6), .GND_b_1_row_4(net1650[0:6]), .Vs_b_0_row_4(net112[0:6]), .Vs_b_1_row_4(net113[0:6]), .VINJ_b_1_row_4(net1656[0:6]), .Vsel_b_0_row_4(net1620[0:6]), .Vsel_b_1_row_4(net1621[0:6]), .Vg_b_0_row_4(net1632[0:6]), .Vg_b_1_row_4(net1633[0:6]), .VTUN_brow_4(net1644[0:6]), .Vd_Rl_0_col_0(net1985[0:5]), .Vd_Rl_1_col_0(net1986[0:5]), .Vd_Rl_2_col_0(net1987[0:5]), .Vd_Rl_3_col_0(net1988[0:5]), .Vd_Pl_0_col_0(net1816[0:5]), .Vd_Pl_1_col_0(net1817[0:5]), .Vd_Pl_2_col_0(net1818[0:5]), .Vd_Pl_3_col_0(net1819[0:5]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(6), .GND_b_1_row_4(net1689[0:6]), .Vs_b_0_row_4(net237[0:6]), .Vs_b_1_row_4(net236[0:6]), .VINJ_b_1_row_4(net1688[0:6]), .Vsel_b_0_row_4(net1690[0:6]), .Vsel_b_1_row_4(net1692[0:6]), .Vg_b_0_row_4(net1691[0:6]), .Vg_b_1_row_4(net1693[0:6]), .VTUN_brow_4(net1687[0:6]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(22), .matrix_row(5), .matrix_col(1), .A_0_col_0(net2019[0:5]), .A_1_col_0(net2020[0:5]), .A_2_col_0(net2021[0:5]), .A_3_col_0(net2022[0:5]), .Prog_brow_4(net1978[0:1]), .VDD_brow_4(net1957[0:1]), .GND_brow_4(net1689[5:6]), .Progrow_0(net1978[0:1]));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(6), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1666[0:1]), .Vsel_b_0_row_4(net1669[0:1]), .Vsel_b_1_row_4(net1670[0:1]), .Vg_b_0_row_4(net1671[0:1]), .Vg_b_1_row_4(net1672[0:1]), .VTUN_brow_4(net1667[0:1]), .GND_b_1_row_4(net1668[0:1]));
	S_BLOCK_BUFFER I__4 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__5 (.island_num(0), .row(0), .col(8), .matrix_row(4), .matrix_col(1), .n_0_row_0(net1926[0:1]), .n_1_row_0(net1927[0:1]), .n_2_row_0(net1928[0:1]), .n_3_row_0(net1929[0:1]));
	S_BLOCK_CONN_PINS I__6 (.island_num(0), .row(4), .col(8), .matrix_row(1), .matrix_col(1), .s_0_row_0(net1958), .s_1_row_0(net1959), .s_2_row_0(net1960), .s_3_row_0(net1961));
	S_BLOCK_SPACE_UP_PINS I__7 (.island_num(0), .row(0), .col(9), .matrix_row(3), .matrix_col(1), .n_0_row_0(net1930[0:1]), .n_1_row_0(net1931[0:1]), .n_2_row_0(net1932[0:1]), .n_3_row_0(net1933[0:1]));
	S_BLOCK_CONN_PINS I__8 (.island_num(0), .row(3), .col(9), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__9 (.island_num(0), .row(4), .col(9), .matrix_row(1), .matrix_col(1), .s_0_row_0(net1962), .s_1_row_0(net1963), .s_2_row_0(net1964), .s_3_row_0(net1965));
	S_BLOCK_SPACE_UP_PINS I__10 (.island_num(0), .row(0), .col(10), .matrix_row(2), .matrix_col(1), .n_0_row_0(net1934[0:1]), .n_1_row_0(net1935[0:1]), .n_2_row_0(net1936[0:1]), .n_3_row_0(net1937[0:1]));
	S_BLOCK_CONN_PINS I__11 (.island_num(0), .row(2), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__12 (.island_num(0), .row(3), .col(10), .matrix_row(2), .matrix_col(1), .s_0_row_1(net1966[0:1]), .s_1_row_1(net1967[0:1]), .s_2_row_1(net1968[0:1]), .s_3_row_1(net1969[0:1]));
	S_BLOCK_SPACE_UP_PINS I__13 (.island_num(0), .row(0), .col(11), .matrix_row(1), .matrix_col(1), .n_0_row_0(net1938), .n_1_row_0(net1939), .n_2_row_0(net1940), .n_3_row_0(net1941));
	S_BLOCK_CONN_PINS I__14 (.island_num(0), .row(1), .col(11), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__15 (.island_num(0), .row(2), .col(11), .matrix_row(3), .matrix_col(1), .s_0_row_2(net1970[0:1]), .s_1_row_2(net1971[0:1]), .s_2_row_2(net1972[0:1]), .s_3_row_2(net1973[0:1]));
	S_BLOCK_CONN_PINS I__16 (.island_num(0), .row(0), .col(12), .matrix_row(1), .matrix_col(1), .n_0_row_0(net1942), .n_1_row_0(net1943), .n_2_row_0(net1944), .n_3_row_0(net1945));
	S_BLOCK_SPACE_DOWN_PINS I__17 (.island_num(0), .row(1), .col(12), .matrix_row(4), .matrix_col(1), .s_0_row_3(net1974[0:1]), .s_1_row_3(net1975[0:1]), .s_2_row_3(net1976[0:1]), .s_3_row_3(net1977[0:1]));
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(13), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1673[0:1]), .Vsel_b_0_row_4(net1676[0:1]), .Vsel_b_1_row_4(net1677[0:1]), .Vg_b_0_row_4(net1678[0:1]), .Vg_b_1_row_4(net1679[0:1]), .VTUN_brow_4(net1674[0:1]), .GND_b_1_row_4(net1675[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1680[0:1]), .Vsel_b_0_row_4(net1683[0:1]), .Vsel_b_1_row_4(net1684[0:1]), .Vg_b_0_row_4(net1685[0:1]), .Vg_b_1_row_4(net1686[0:1]), .VTUN_brow_4(net1681[0:1]), .GND_b_1_row_4(net1682[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(5), .decode_n1_VGRUN_2_(net1922[0]), .decode_n1_VGRUN_3_(net1923[0]), .decode_n2_VGRUN_0_(net1924[0]), .decode_n2_VGRUN_1_(net1925[0]), .decode_n5_VGRUN_2_(net2005[0]), .decode_n5_VGRUN_3_(net2006[0]), .decode_n6_VGRUN_0_(net2007[0]), .decode_n6_VGRUN_1_(net2008[0]), .decode_n4_n0_RUN_OUT_0_(net1792[0]), .decode_n4_n0_RUN_OUT_1_(net1793[0]), .decode_n4_n0_RUN_OUT_2_(net1794[0]), .decode_n4_n0_RUN_OUT_3_(net1795[0]), .decode_n4_n1_RUN_OUT_0_(net1796[0]), .decode_n4_n1_RUN_OUT_1_(net1797[0]), .decode_n4_n1_RUN_OUT_2_(net1784), .decode_n4_n1_RUN_OUT_3_(net1785), .decode_n4_n2_RUN_OUT_0_(net1786), .decode_n4_n2_RUN_OUT_1_(net1787), .decode_n4_n2_RUN_OUT_2_(net1798[0]), .decode_n4_n2_RUN_OUT_3_(net1799[0]), .decode_n4_n3_RUN_OUT_0_(net1800[0]), .decode_n4_n3_RUN_OUT_1_(net1801[0]), .decode_n4_n3_RUN_OUT_2_(net1802[0]), .decode_n4_n3_RUN_OUT_3_(net1803[0]), .decode_n4_n4_RUN_OUT_0_(net1804[0]), .decode_n4_n4_RUN_OUT_1_(net1805[0]), .decode_n4_n4_RUN_OUT_2_(net1806[0]), .decode_n4_n4_RUN_OUT_3_(net1807[0]), .decode_n4_n5_RUN_OUT_0_(net1808[0]), .decode_n4_n5_RUN_OUT_1_(net1809[0]), .decode_n4_n5_RUN_OUT_2_(net1788), .decode_n4_n5_RUN_OUT_3_(net1789), .decode_n4_n6_RUN_OUT_0_(net1790), .decode_n4_n6_RUN_OUT_1_(net1791), .decode_n4_n6_RUN_OUT_2_(net1810[0]), .decode_n4_n6_RUN_OUT_3_(net1811[0]), .decode_n4_n7_RUN_OUT_0_(net1812[0]), .decode_n4_n7_RUN_OUT_1_(net1813[0]), .decode_n4_n7_RUN_OUT_2_(net1814[0]), .decode_n4_n7_RUN_OUT_3_(net1815[0]), .decode_n4_n0_OUT_0_(net1730), .decode_n4_n0_OUT_1_(net1731), .decode_n4_n0_OUT_2_(net1734), .decode_n4_n0_OUT_3_(net1735), .decode_n4_n1_OUT_0_(net1738), .decode_n4_n1_OUT_1_(net1739), .decode_n4_n1_OUT_2_(net1742), .decode_n4_n1_OUT_3_(net1743), .decode_n4_n2_OUT_0_(net1746), .decode_n4_n2_OUT_1_(net1747), .decode_n4_n2_OUT_2_(net1750), .decode_n4_n2_OUT_3_(net1751), .decode_n4_n3_OUT_0_(net1754), .decode_n4_n3_OUT_1_(net1755), .decode_n4_n4_OUT_0_(net1758), .decode_n4_n4_OUT_1_(net1759), .decode_n4_n4_OUT_2_(net1762), .decode_n4_n4_OUT_3_(net1763), .decode_n4_n5_OUT_0_(net1766), .decode_n4_n5_OUT_1_(net1767), .decode_n4_n5_OUT_2_(net1770), .decode_n4_n5_OUT_3_(net1771), .decode_n4_n6_OUT_0_(net1774), .decode_n4_n6_OUT_1_(net1775), .decode_n4_n6_OUT_2_(net1778), .decode_n4_n6_OUT_3_(net1779), .decode_n4_n7_OUT_0_(net1782), .decode_n4_n7_OUT_1_(net1783), .decode_n0_ENABLE(net1946), .decode_n4_n0_VINJ_b_0_(net1728), .decode_n4_n0_VINJ_b_1_(net1732), .decode_n4_n1_VINJ_b_0_(net1736), .decode_n4_n1_VINJ_b_1_(net1740), .decode_n4_n2_VINJ_b_0_(net1744), .decode_n4_n2_VINJ_b_1_(net1748), .decode_n4_n3_VINJ_b_0_(net1752), .decode_n4_n4_VINJ_b_0_(net1756), .decode_n4_n4_VINJ_b_1_(net1760), .decode_n4_n5_VINJ_b_0_(net1764), .decode_n4_n5_VINJ_b_1_(net1768), .decode_n4_n6_VINJ_b_0_(net1772), .decode_n4_n6_VINJ_b_1_(net1776), .decode_n4_n7_VINJ_b_0_(net1780), .decode_n4_n0_GND_b_0_(net1729), .decode_n4_n0_GND_b_1_(net1733), .decode_n4_n1_GND_b_0_(net1737), .decode_n4_n1_GND_b_1_(net1741), .decode_n4_n2_GND_b_0_(net1745), .decode_n4_n2_GND_b_1_(net1749), .decode_n4_n3_GND_b_0_(net1753), .decode_n4_n4_GND_b_0_(net1757), .decode_n4_n4_GND_b_1_(net1761), .decode_n4_n5_GND_b_0_(net1765), .decode_n4_n5_GND_b_1_(net1769), .decode_n4_n6_GND_b_0_(net1773), .decode_n4_n6_GND_b_1_(net1777), .decode_n4_n7_GND_b_0_(net1781), .decode_n0_VINJV(net1953), .decode_n0_GNDV(net1955));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(22), .switch_n3_VPWR_0_(net1784), .switch_n3_VPWR_1_(net1785), .switch_n4_VPWR_0_(net1786), .switch_n4_VPWR_1_(net1787), .switch_n17_VPWR_0_(net1788), .switch_n17_VPWR_1_(net1789), .switch_n18_VPWR_0_(net1790), .switch_n18_VPWR_1_(net1791), .switch_n0_RUN_IN_0_(net1921), .switch_n0_RUN_IN_1_(net1921), .switch_n1_RUN_IN_0_(net1921), .switch_n1_RUN_IN_1_(net1921), .switch_n2_RUN_IN_0_(net1921), .switch_n2_RUN_IN_1_(net1921), .switch_n3_RUN_IN_0_(net1921), .switch_n3_RUN_IN_1_(net1921), .switch_n4_RUN_IN_0_(net1921), .switch_n4_RUN_IN_1_(net1921), .switch_n5_RUN_IN_0_(net1921), .switch_n5_RUN_IN_1_(net1921), .switch_n6_RUN_IN_0_(net1921), .switch_n6_RUN_IN_1_(net1921), .switch_n13_RUN_IN_0_(net1921), .switch_n13_RUN_IN_1_(net1921), .switch_n15_RUN_IN_0_(net1921), .switch_n15_RUN_IN_1_(net1921), .switch_n16_RUN_IN_0_(net1921), .switch_n16_RUN_IN_1_(net1921), .switch_n17_RUN_IN_0_(net1921), .switch_n17_RUN_IN_1_(net1921), .switch_n18_RUN_IN_0_(net1921), .switch_n18_RUN_IN_1_(net1921), .switch_n19_RUN_IN_0_(net1921), .switch_n19_RUN_IN_1_(net1921), .switch_n20_RUN_IN_0_(net1921), .switch_n20_RUN_IN_1_(net1921), .switch_n21_RUN_IN_0_(net1921), .switch_n21_RUN_IN_1_(net1921), .switch_n0_GND_T(net1729), .switch_n1_GND_T(net1733), .switch_n2_GND_T(net1737), .switch_n3_GND_T(net1741), .switch_n4_GND_T(net1745), .switch_n5_GND_T(net1749), .switch_n6_GND_T(net1753), .switch_n14_GND_T(net1757), .switch_n15_GND_T(net1761), .switch_n16_GND_T(net1765), .switch_n17_GND_T(net1769), .switch_n18_GND_T(net1773), .switch_n19_GND_T(net1777), .switch_n20_GND_T(net1781), .switch_n0_VTUN_T(net2010[0]), .switch_n0_decode_0_(net1730), .switch_n0_decode_1_(net1731), .switch_n1_decode_0_(net1734), .switch_n1_decode_1_(net1735), .switch_n2_decode_0_(net1738), .switch_n2_decode_1_(net1739), .switch_n3_decode_0_(net1742), .switch_n3_decode_1_(net1743), .switch_n4_decode_0_(net1746), .switch_n4_decode_1_(net1747), .switch_n5_decode_0_(net1750), .switch_n5_decode_1_(net1751), .switch_n6_decode_0_(net1754), .switch_n6_decode_1_(net1755), .switch_n14_decode_0_(net1758), .switch_n14_decode_1_(net1759), .switch_n15_decode_0_(net1762), .switch_n15_decode_1_(net1763), .switch_n16_decode_0_(net1766), .switch_n16_decode_1_(net1767), .switch_n17_decode_0_(net1770), .switch_n17_decode_1_(net1771), .switch_n18_decode_0_(net1774), .switch_n18_decode_1_(net1775), .switch_n19_decode_0_(net1778), .switch_n19_decode_1_(net1779), .switch_n20_decode_0_(net1782), .switch_n20_decode_1_(net1783), .switch_n0_VINJ_T(net1728), .switch_n1_VINJ_T(net1732), .switch_n2_VINJ_T(net1736), .switch_n3_VINJ_T(net1740), .switch_n4_VINJ_T(net1744), .switch_n5_VINJ_T(net1748), .switch_n6_VINJ_T(net1752), .switch_n14_VINJ_T(net1756), .switch_n15_VINJ_T(net1760), .switch_n16_VINJ_T(net1764), .switch_n17_VINJ_T(net1768), .switch_n18_VINJ_T(net1772), .switch_n19_VINJ_T(net1776), .switch_n20_VINJ_T(net1780), .switch_n0_RUN(net1979), .switch_n0_vgsel_r(net1980));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5), .decode_n0_IN_0_(net2018), .decode_n0_IN_1_(net2017), .decode_n0_IN_2_(net2016), .decode_n0_IN_3_(net2015), .decode_n0_IN_4_(net2014), .decode_n0_ENABLE(net2044));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select), .switch_n0_prog_drainrail(net1947), .switch_n0_run_drainrail(net1948), .switch_n0_VINJ(net1954), .switch_n0_GND(net1956));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch), .switch_n0_PR_0_(net1816[0]), .switch_n0_PR_1_(net1817[0]), .switch_n0_PR_2_(net1818[0]), .switch_n0_PR_3_(net1819[0]), .switch_n1_PR_0_(net1816[1]), .switch_n1_PR_1_(net1817[1]), .switch_n1_PR_2_(net1818[1]), .switch_n1_PR_3_(net1819[1]), .switch_n2_PR_0_(net1816[2]), .switch_n2_PR_1_(net1817[2]), .switch_n2_PR_2_(net1818[2]), .switch_n2_PR_3_(net1819[2]), .switch_n3_PR_0_(net1816[3]), .switch_n3_PR_1_(net1817[3]), .switch_n3_PR_2_(net1818[3]), .switch_n3_PR_3_(net1819[3]), .switch_n4_PR_0_(net1816[4]), .switch_n4_PR_1_(net1817[4]), .switch_n4_PR_2_(net1818[4]), .switch_n4_PR_3_(net1819[4]), .switch_n0_In_0_(net1985[0]), .switch_n0_In_1_(net1986[0]), .switch_n0_In_2_(net1987[0]), .switch_n0_In_3_(net1988[0]), .switch_n1_In_0_(net1985[1]), .switch_n1_In_1_(net1986[1]), .switch_n1_In_2_(net1987[1]), .switch_n1_In_3_(net1988[1]), .switch_n2_In_0_(net1985[2]), .switch_n2_In_1_(net1986[2]), .switch_n2_In_2_(net1987[2]), .switch_n2_In_3_(net1988[2]), .switch_n3_In_0_(net1985[3]), .switch_n3_In_1_(net1986[3]), .switch_n3_In_2_(net1987[3]), .switch_n3_In_3_(net1988[3]), .switch_n4_In_0_(net1985[4]), .switch_n4_In_1_(net1986[4]), .switch_n4_In_2_(net1987[4]), .switch_n4_In_3_(net1988[4]), .switch_n0_VDD(net1954), .switch_n0_GND(net1956), .switch_n0_RUN(net1979));
	none switch_ind(.island_num(0), .direction(horizontal), .col(7));
	none switch_ind(.island_num(0), .direction(horizontal), .col(8));
	none switch_ind(.island_num(0), .direction(horizontal), .col(9));
	none switch_ind(.island_num(0), .direction(horizontal), .col(10));
	none switch_ind(.island_num(0), .direction(horizontal), .col(11));
	none switch_ind(.island_num(0), .direction(horizontal), .col(12));
	none switch_ind(.island_num(0), .direction(horizontal), .col(14));


	/* Island 1 */
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__0 (.island_num(1), .row(0), .col(0), .matrix_row(1), .matrix_col(7));
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(5), .matrix_col(7), .GND_b_0_row_4(net882[0:7]), .GND_b_1_row_4(net883[0:7]), .Vs_b_0_row_4(net890[0:7]), .Vs_b_1_row_4(net891[0:7]), .VINJ_b_0_row_4(net892[0:7]), .VINJ_b_1_row_4(net893[0:7]), .Vsel_b_0_row_4(net894[0:7]), .Vsel_b_1_row_4(net895[0:7]), .Vg_b_0_row_4(net896[0:7]), .Vg_b_1_row_4(net897[0:7]), .VTUN_brow_4(net898[0:7]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(7), .matrix_row(1), .matrix_col(7));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(7), .matrix_row(4), .matrix_col(7));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(5), .col(7), .matrix_row(1), .matrix_col(7));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(14), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1546), .P_1_row_0(net1547), .A_0_row_0(net1548), .A_1_row_0(net1549), .A_2_row_0(net1550), .A_3_row_0(net1551), .Progrow_0(net1917), .VDDrow_0(net1957[0]), .GNDrow_0(net1689[5]));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(14), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1561), .P_1_row_0(net1562), .A_0_row_0(net1563), .A_1_row_0(net1564), .A_2_row_0(net1565), .A_3_row_0(net1566));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(14), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1579), .P_1_row_0(net1580), .P_2_row_0(net1581), .P_3_row_0(net1582), .A_0_row_0(net1583), .A_1_row_0(net1584));
	TSMC350nm_4TGate_ST_BMatrix_NoSwitch I__8 (.island_num(1), .row(3), .col(14), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1594), .P_1_row_0(net1595), .P_2_row_0(net1596), .P_3_row_0(net1597), .A_0_row_0(net1598), .A_1_row_0(net1599), .A_2_row_0(net1600), .A_3_row_0(net1601));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(14), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1613), .A_1_row_0(net1614), .A_2_row_0(net1615), .A_3_row_0(net1616));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(14), .matrix_row(1), .matrix_col(1), .Prog_brow_0(net1920[0]), .VDD_brow_0(net1919[0]), .GND_brow_0(net1918[0]));
	TSMC350nm_OutMtrx_IndrctSwcs I__11 (.island_num(1), .row(7), .col(7), .matrix_row(1), .matrix_col(7));
	TSMC350nm_4x2_Indirect I__12 (.island_num(1), .row(8), .col(7), .matrix_row(2), .matrix_col(7), .Vd_Rl_0_col_0(net1403[0:2]), .Vd_Rl_1_col_0(net1404[0:2]), .Vd_Rl_2_col_0(net1405[0:2]), .Vd_Rl_3_col_0(net1406[0:2]), .Vd_Pl_0_col_0(net1407[0:2]), .Vd_Pl_1_col_0(net1408[0:2]), .Vd_Pl_2_col_0(net1409[0:2]), .Vd_Pl_3_col_0(net1410[0:2]));
	TSMC350nm_4TGate_ST_BMatrix I__13 (.island_num(1), .row(8), .col(14), .matrix_row(2), .matrix_col(1), .A_0_col_0(net1949[0:2]), .A_1_col_0(net1950[0:2]), .A_2_col_0(net1951[0:2]), .A_3_col_0(net1952[0:2]), .Progrow_0(net1920[0:1]), .VDDrow_0(net1919[0:1]), .GNDrow_0(net1918[0:1]));
	TSMC350nm_TA2Cell_Weak cab_device_14 (.island_num(1), .row(2), .col(15), .VD_P_0_(net1546), .VD_P_1_(net1547), .VIN1_PLUS(net1548), .VIN1_MINUS(net1549), .VIN2_PLUS(net1550), .VIN2_MINUS(net1551), .OUTPUT_0_(net1552[0]), .OUTPUT_1_(net1553[0]), .Vsel_0_(net1608), .Vsel_1_(net1554), .RUN(net1555), .Vg_0_(net1556), .Vg_1_(net1557), .PROG(net1978[0]), .VTUN(net1558), .VINJ(net1559), .GND(net1560), .VPWR(net2013[0]), .Vsel_b_0_(net1569), .Vsel_b_1_(net1570), .RUN_b(net1571), .Vg_b_0_(net1572), .Vg_b_1_(net1573), .PROG_b(net1574), .VTUN_b(net1575), .VINJ_b(net1576), .GND_b(net1577), .VPWR_b(net1578));
	TSMC350nm_TA2Cell_Strong cab_device_15 (.island_num(1), .row(3), .col(15), .VD_P_0_(net1561), .VD_P_1_(net1562), .VIN1_PLUS(net1563), .VIN1_MINUS(net1564), .VIN2_PLUS(net1565), .VIN2_MINUS(net1566), .OUTPUT_0_(net1567[0]), .OUTPUT_1_(net1568[0]), .Vsel_0_(net1569), .Vsel_1_(net1570), .RUN(net1571), .Vg_0_(net1572), .Vg_1_(net1573), .PROG(net1574), .VTUN(net1575), .VINJ(net1576), .GND(net1577), .VPWR(net1578), .Vsel_b_0_(net1588), .Vsel_b_1_(net1589), .Vg_b_0_(net1590), .Vg_b_1_(net1591), .VTUN_b(net1593), .VINJ_b(net1587), .GND_b(net1592));
	TSMC350nm_Cap_Bank cab_device_16 (.island_num(1), .row(4), .col(15), .VD_P_0_(net1579), .VD_P_1_(net1580), .VD_P_2_(net1581), .VD_P_3_(net1582), .VIN_0_(net1583), .VIN_1_(net1584), .OUT_0_(net1585[0]), .OUT_1_(net1586[0]), .VINJ(net1587), .Vsel_0_(net1588), .Vsel_1_(net1589), .Vg_0_(net1590), .Vg_1_(net1591), .GND(net1592), .VTUN(net1593), .VINJ_b(net1609), .Vg_b_0_(net1610), .GND_b(net1612), .VTUN_b(net1611));
	TSMC350nm_4WTA_IndirectProg cab_device_17 (.island_num(1), .row(5), .col(15), .VD_P_0_(net1594), .VD_P_1_(net1595), .VD_P_2_(net1596), .VD_P_3_(net1597), .Iin_0_(net1598), .Iin_1_(net1599), .Iin_2_(net1600), .Iin_3_(net1601), .Vout_0_(net1602[0]), .Vout_1_(net1603[0]), .Vout_2_(net1604[0]), .Vout_3_(net1605[0]), .Vmid(net1606[0]), .Vbias(net1607[0]), .Vsel(net1608), .Vs(net2013[0]), .VINJ(net1609), .Vg(net1610), .VTUN(net1611), .GND(net1612), .PROG(net1978[0]), .GND_b(net1619));
	TSMC350nm_NandPfets cab_device_18 (.island_num(1), .row(6), .col(15), .GATE_N(net1613), .SOURCE_N(net1614), .GATE_P(net1615), .SOURCE_P(net1616), .DRAIN_N(net1617[0]), .DRAIN_P(net1618[0]), .VPWR(net2013[0]), .GND(net1619));
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6), .decode_n0_IN_0_(net2043), .decode_n0_IN_1_(net2042), .decode_n0_IN_2_(net2041), .decode_n0_IN_3_(net2040), .decode_n0_IN_4_(net2039), .decode_n0_ENABLE(net2044));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(1), .direction(vertical), .num(10), .type(drain_select), .switch_n0_prog_drainrail(net1947), .switch_n0_run_drainrail(net1948));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(10), .type(prog_switch), .switch_n6_PR_0_(net1901[0]), .switch_n6_PR_1_(net1905[0]), .switch_n6_PR_2_(net1909[0]), .switch_n6_PR_3_(net1913[0]), .switch_n6_In_0_(net1900[0]), .switch_n6_In_1_(net1904[0]), .switch_n6_In_2_(net1908[0]), .switch_n6_In_3_(net1912[0]), .switch_n0_RUN(net1979));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(16), .switch_n0_Input_0_(net1957[0]), .switch_n0_Input_1_(net1650[0]), .switch_n1_Input_0_(net112[1]), .switch_n1_Input_1_(net113[1]), .switch_n2_Input_0_(net112[2]), .switch_n2_Input_1_(net113[2]), .switch_n3_Input_0_(net237[0]), .switch_n6_Input_1_(net1899[0]), .switch_n7_Input_0_(net1552[0]), .switch_n7_Input_1_(net1553[0]), .switch_n8_Input_0_(net1567[0]), .switch_n8_Input_1_(net1568[0]), .switch_n9_Input_0_(net1585[0]), .switch_n9_Input_1_(net1586[0]), .switch_n10_Input_0_(net1602[0]), .switch_n10_Input_1_(net1603[0]), .switch_n11_Input_0_(net1604[0]), .switch_n11_Input_1_(net1605[0]), .switch_n12_Input_0_(net1606[0]), .switch_n12_Input_1_(net1607[0]), .switch_n13_Input_0_(net1617[0]), .switch_n13_Input_1_(net1618[0]), .switch_n0_GND(net1650[0]), .switch_n1_GND(net1650[1]), .switch_n2_GND(net1650[2]), .switch_n3_GND(net1650[3]), .switch_n4_GND(net1650[4]), .switch_n5_GND(net1650[5]), .switch_n6_GND(net1668[0]), .switch_n7_GND(net1675[0]), .switch_n8_GND(net1682[0]), .switch_n9_GND(net1689[0]), .switch_n10_GND(net1689[1]), .switch_n11_GND(net1689[2]), .switch_n12_GND(net1689[3]), .switch_n13_GND(net1689[4]), .switch_n14_GND(net1689[5]), .switch_n0_Vsel_0_(net1620[0]), .switch_n0_Vsel_1_(net1621[0]), .switch_n1_Vsel_0_(net1620[1]), .switch_n1_Vsel_1_(net1621[1]), .switch_n2_Vsel_0_(net1620[2]), .switch_n2_Vsel_1_(net1621[2]), .switch_n3_Vsel_0_(net1620[3]), .switch_n3_Vsel_1_(net1621[3]), .switch_n4_Vsel_0_(net1620[4]), .switch_n4_Vsel_1_(net1621[4]), .switch_n5_Vsel_0_(net1620[5]), .switch_n5_Vsel_1_(net1621[5]), .switch_n6_Vsel_0_(net1670[0]), .switch_n6_Vsel_1_(net1669[0]), .switch_n7_Vsel_0_(net1677[0]), .switch_n7_Vsel_1_(net1676[0]), .switch_n8_Vsel_0_(net1684[0]), .switch_n8_Vsel_1_(net1683[0]), .switch_n9_Vsel_0_(net1690[0]), .switch_n9_Vsel_1_(net1692[0]), .switch_n10_Vsel_0_(net1690[1]), .switch_n10_Vsel_1_(net1692[1]), .switch_n11_Vsel_0_(net1690[2]), .switch_n11_Vsel_1_(net1692[2]), .switch_n12_Vsel_0_(net1690[3]), .switch_n12_Vsel_1_(net1692[3]), .switch_n13_Vsel_0_(net1690[4]), .switch_n13_Vsel_1_(net1692[4]), .switch_n14_Vsel_0_(net1690[5]), .switch_n14_Vsel_1_(net1692[5]), .switch_n0_Vg_global_0_(net1632[0]), .switch_n0_Vg_global_1_(net1633[0]), .switch_n1_Vg_global_0_(net1632[1]), .switch_n1_Vg_global_1_(net1633[1]), .switch_n2_Vg_global_0_(net1632[2]), .switch_n2_Vg_global_1_(net1633[2]), .switch_n3_Vg_global_0_(net1632[3]), .switch_n3_Vg_global_1_(net1633[3]), .switch_n4_Vg_global_0_(net1632[4]), .switch_n4_Vg_global_1_(net1633[4]), .switch_n5_Vg_global_0_(net1632[5]), .switch_n5_Vg_global_1_(net1633[5]), .switch_n6_Vg_global_0_(net1672[0]), .switch_n6_Vg_global_1_(net1671[0]), .switch_n7_Vg_global_0_(net1679[0]), .switch_n7_Vg_global_1_(net1678[0]), .switch_n8_Vg_global_0_(net1686[0]), .switch_n8_Vg_global_1_(net1685[0]), .switch_n9_Vg_global_0_(net1691[0]), .switch_n9_Vg_global_1_(net1693[0]), .switch_n10_Vg_global_0_(net1691[1]), .switch_n10_Vg_global_1_(net1693[1]), .switch_n11_Vg_global_0_(net1691[2]), .switch_n11_Vg_global_1_(net1693[2]), .switch_n12_Vg_global_0_(net1691[3]), .switch_n12_Vg_global_1_(net1693[3]), .switch_n13_Vg_global_0_(net1691[4]), .switch_n13_Vg_global_1_(net1693[4]), .switch_n14_Vg_global_0_(net1691[5]), .switch_n14_Vg_global_1_(net1693[5]), .switch_n0_VTUN(net1644[0]), .switch_n1_VTUN(net1644[1]), .switch_n2_VTUN(net1644[2]), .switch_n3_VTUN(net1644[3]), .switch_n4_VTUN(net1644[4]), .switch_n5_VTUN(net1644[5]), .switch_n6_VTUN(net1667[0]), .switch_n7_VTUN(net1674[0]), .switch_n8_VTUN(net1681[0]), .switch_n9_VTUN(net1687[0]), .switch_n10_VTUN(net1687[1]), .switch_n11_VTUN(net1687[2]), .switch_n12_VTUN(net1687[3]), .switch_n13_VTUN(net1687[4]), .switch_n14_VTUN(net1687[5]), .switch_n0_VINJ(net1656[0]), .switch_n1_VINJ(net1656[1]), .switch_n2_VINJ(net1656[2]), .switch_n3_VINJ(net1656[3]), .switch_n4_VINJ(net1656[4]), .switch_n5_VINJ(net1656[5]), .switch_n6_VINJ(net1666[0]), .switch_n7_VINJ(net1673[0]), .switch_n8_VINJ(net1680[0]), .switch_n9_VINJ(net1688[0]), .switch_n10_VINJ(net1688[1]), .switch_n11_VINJ(net1688[2]), .switch_n12_VINJ(net1688[3]), .switch_n13_VINJ(net1688[4]), .switch_n14_VINJ(net1688[5]), .switch_n0_Vgrun_r(net2009), .switch_n0_Vgrun(net1921), .switch_n0_AVDD_r(net2013[0]), .switch_n0_run_r(net1916), .switch_n0_prog_r(net1917), .switch_n0_run(net1979));
	none switch_ind(.island_num(1), .direction(horizontal), .col(14));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(15), .VPWR_0_(net1957[0]), .VPWR_1_(net1957[0]), .RUN_IN_0_(net2009), .RUN_IN_1_(net2009), .GND_T(net1689[5]), .VTUN_T(net1687[5]), .decode_0_(net1690[5]), .decode_1_(net1692[5]), .VINJ_T(net1688[5]), .GND(net1560), .CTRL_B_0_(net1608), .CTRL_B_1_(net1554), .run_r(net1555), .prog_r(net1978[0]), .Vg_0_(net1556), .Vg_1_(net1557), .VTUN(net1558), .VINJ(net1559), .VDD_1_(net2013[0]), .PROG(net1917), .RUN(net1916), .Vgsel(net1980));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net890[0:6]), .out_1_row_0(net891[0:6]), .VINJ_0_row_0(net892[0:6]), .VINJ_1_row_0(net893[0:6]), .Vsel_0_row_0(net894[0:6]), .Vsel_1_row_0(net895[0:6]), .Vg_0_row_0(net896[0:6]), .Vg_1_row_0(net897[0:6]), .GNDrow_0(net882[0:6]), .VTUNrow_0(net898[0:6]), .Dcol_0(net112[5:6]), .CLKcol_0(net113[5:6]), .Qcol_5(net236[3:4]), .comcol_0(net1899[0:1]), .VDDcol_0(net2013[0:1]), .Vd_Pcol_0(net1913[0:1]), .Vd_in_0_col_0(net1900[0:1]), .Vd_in_1_col_0(net1904[0:1]), .Vd_in_2_col_0(net1908[0:1]), .Vd_in_3_col_0(net1912[0:1]), .Vd_in_4_col_0(net1901[0:1]), .Vd_in_5_col_0(net1905[0:1]), .Vd_in_6_col_0(net1909[0:1]), .Vd_in_7_col_0(net1913[0:1]), .Vd_o_0_col_5(net1403[0:1]), .Vd_o_1_col_5(net1404[0:1]), .Vd_o_2_col_5(net1405[0:1]), .Vd_o_3_col_5(net1406[0:1]), .Vd_o_4_col_5(net1407[0:1]), .Vd_o_5_col_5(net1408[0:1]), .Vd_o_6_col_5(net1409[0:1]), .Vd_o_7_col_5(net1410[0:1]));

 	/*Programming Mux */ 


	/* Frame */ 
	tile_analog_frame cab_frame(.pin_layer(METAL3), .N_n_gateEN(net1946), .N_n_programdrain(net1947), .N_n_rundrain(net1948), .N_n_cew0(net1922[0]), .N_n_cew1(net1923[0]), .N_n_cew2(net1924[0]), .N_n_cew3(net1925[0]), .N_n_vtun(net2010[0]), .N_n_vinj_0_(net1953), .N_n_vinj_1_(net1954), .N_n_vinj_2_(net1688[5]), .N_n_gnd_0_(net1955), .N_n_gnd_1_(net1956), .N_n_gnd_2_(net1689[5]), .N_n_avdd(net1957[0]), .N_n_s0(net1926[0]), .N_n_s1(net1927[0]), .N_n_s2(net1928[0]), .N_n_s3(net1929[0]), .N_n_s4(net1930[0]), .N_n_s5(net1931[0]), .N_n_s6(net1932[0]), .N_n_s7(net1933[0]), .N_n_s8(net1934[0]), .N_n_s9(net1935[0]), .N_n_s10(net1936[0]), .N_n_s11(net1937[0]), .N_n_s12(net1938), .N_n_s13(net1939), .N_n_s14(net1940), .N_n_s15(net1941), .N_n_s16(net1942), .N_n_s17(net1943), .N_n_s18(net1944), .N_n_s19(net1945), .N_n_prog(net1978[0]), .N_n_run(net1979), .N_n_vgsel(net1980), .S_s_gateEN(net1946), .S_s_programdrain(net1947), .S_s_rundrain(net1948), .S_s_cew0(net1949[0]), .S_s_cew1(net1950[0]), .S_s_cew2(net1951[0]), .S_s_cew3(net1952[0]), .S_s_vtun(net2010[0]), .S_s_vinj_0_(net1953), .S_s_vinj_1_(net1954), .S_s_vinj_2_(net1688[5]), .S_s_gnd_0_(net1955), .S_s_gnd_1_(net1956), .S_s_gnd_2_(net1689[5]), .S_s_avdd(net1957[0]), .S_s_s0(net1958), .S_s_s1(net1959), .S_s_s2(net1960), .S_s_s3(net1961), .S_s_s4(net1962), .S_s_s5(net1963), .S_s_s6(net1964), .S_s_s7(net1965), .S_s_s8(net1966[0]), .S_s_s9(net1967[0]), .S_s_s10(net1968[0]), .S_s_s11(net1969[0]), .S_s_s12(net1970[0]), .S_s_s13(net1971[0]), .S_s_s14(net1972[0]), .S_s_s15(net1973[0]), .S_s_s16(net1974[0]), .S_s_s17(net1975[0]), .S_s_s18(net1976[0]), .S_s_s19(net1977[0]), .S_s_prog(net1978[0]), .S_s_run(net1979), .S_s_vgsel(net1980), .W_w_cns0(net1949[1]), .W_w_cns1(net1950[1]), .W_w_cns2(net1951[1]), .W_w_cns3(net1952[1]), .W_w_vgrun(net2009), .W_w_vtun(net2010[0]), .W_w_vinj(net1688[5]), .W_w_gnd(net1689[5]), .W_w_avdd(net2013[0]), .W_w_drainbit4(net2014), .W_w_drainbit3(net2015), .W_w_drainbit2(net2016), .W_w_drainbit1(net2017), .W_w_drainbit0(net2018), .W_w_s0(net1985[0]), .W_w_s1(net1986[0]), .W_w_s2(net1987[0]), .W_w_s3(net1988[0]), .W_w_s4(net1985[1]), .W_w_s5(net1986[1]), .W_w_s6(net1987[1]), .W_w_s7(net1988[1]), .W_w_s8(net1985[2]), .W_w_s9(net1986[2]), .W_w_s10(net1987[2]), .W_w_s11(net1988[2]), .W_w_s12(net1985[3]), .W_w_s13(net1986[3]), .W_w_s14(net1987[3]), .W_w_s15(net1988[3]), .W_w_s16(net1985[4]), .W_w_s17(net1986[4]), .W_w_s18(net1987[4]), .W_w_s19(net1988[4]), .W_w_drainbit9(net2039), .W_w_drainbit8(net2040), .W_w_drainbit7(net2041), .W_w_drainbit6(net2042), .W_w_drainbit5(net2043), .W_w_drainEN(net2044), .E_e_cns0(net2005[0]), .E_e_cns1(net2006[0]), .E_e_cns2(net2007[0]), .E_e_cns3(net2008[0]), .E_e_vgrun(net2009), .E_e_vtun(net2010[0]), .E_e_vinj(net1688[5]), .E_e_gnd(net1689[5]), .E_e_avdd(net2013[0]), .E_e_drainbit4(net2014), .E_e_drainbit3(net2015), .E_e_drainbit2(net2016), .E_e_drainbit1(net2017), .E_e_drainbit0(net2018), .E_e_s0(net2019[0]), .E_e_s1(net2020[0]), .E_e_s2(net2021[0]), .E_e_s3(net2022[0]), .E_e_s4(net2019[1]), .E_e_s5(net2020[1]), .E_e_s6(net2021[1]), .E_e_s7(net2022[1]), .E_e_s8(net2019[2]), .E_e_s9(net2020[2]), .E_e_s10(net2021[2]), .E_e_s11(net2022[2]), .E_e_s12(net2019[3]), .E_e_s13(net2020[3]), .E_e_s14(net2021[3]), .E_e_s15(net2022[3]), .E_e_s16(net2019[4]), .E_e_s17(net2020[4]), .E_e_s18(net2021[4]), .E_e_s19(net2022[4]), .E_e_drainbit9(net2039), .E_e_drainbit8(net2040), .E_e_drainbit7(net2041), .E_e_drainbit6(net2042), .E_e_drainbit5(net2043), .E_e_drainEN(net2044));
 endmodule