module TOP(port1);


	/* Island 0 */
	TSMC350nm_TA2Cell_Weak I__0 (.island_num(0), .row(0), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net218[0]), .VD_P_1_row_0(net219[0]), .VIN1_PLUSrow_0(net295), .VIN1_MINUSrow_0(net30), .VIN2_PLUSrow_0(net30), .VIN2_MINUSrow_0(net71), .OUTPUT_0_row_0(net30), .OUTPUT_1_row_0(net30), .Vsel_0_row_0(net293), .Vsel_1_row_0(net294), .RUNrow_0(net321), .Vg_0_row_0(net291), .Vg_1_row_0(net292), .PROGrow_0(net320), .VTUNrow_0(net318), .VINJrow_0(net316), .GNDrow_0(net317), .VPWRrow_0(net319));
	TSMC350nm_TA2Cell_Weak I__1 (.island_num(0), .row(1), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net220[0]), .VD_P_1_row_0(net221[0]), .VIN1_PLUSrow_0(net30), .VIN1_MINUSrow_0(net71), .VIN2_PLUSrow_0(net71), .VIN2_MINUSrow_0(net297), .OUTPUT_0_row_0(net71), .OUTPUT_1_row_0(net297));
	TSMC350nm_TA2Cell_Weak I__2 (.island_num(0), .row(2), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net222[0]), .VD_P_1_row_0(net223[0]), .VIN1_PLUSrow_0(net71), .VIN1_MINUSrow_0(net72), .VIN2_PLUSrow_0(net72), .VIN2_MINUSrow_0(net113), .OUTPUT_0_row_0(net72), .OUTPUT_1_row_0(net72));
	TSMC350nm_TA2Cell_Weak I__3 (.island_num(0), .row(3), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net224[0]), .VD_P_1_row_0(net225[0]), .VIN1_PLUSrow_0(net72), .VIN1_MINUSrow_0(net113), .VIN2_PLUSrow_0(net113), .VIN2_MINUSrow_0(net298), .OUTPUT_0_row_0(net113), .OUTPUT_1_row_0(net298));
	TSMC350nm_TA2Cell_Weak I__4 (.island_num(0), .row(4), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net226[0]), .VD_P_1_row_0(net227[0]), .VIN1_PLUSrow_0(net113), .VIN1_MINUSrow_0(net114), .VIN2_PLUSrow_0(net114), .VIN2_MINUSrow_0(net155), .OUTPUT_0_row_0(net114), .OUTPUT_1_row_0(net114));
	TSMC350nm_TA2Cell_Weak I__5 (.island_num(0), .row(5), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net228[0]), .VD_P_1_row_0(net229[0]), .VIN1_PLUSrow_0(net114), .VIN1_MINUSrow_0(net155), .VIN2_PLUSrow_0(net155), .VIN2_MINUSrow_0(net299), .OUTPUT_0_row_0(net155), .OUTPUT_1_row_0(net299));
	TSMC350nm_TA2Cell_Weak I__6 (.island_num(0), .row(6), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net230[0]), .VD_P_1_row_0(net231[0]), .VIN1_PLUSrow_0(net155), .VIN1_MINUSrow_0(net156), .VIN2_PLUSrow_0(net156), .VIN2_MINUSrow_0(net195), .OUTPUT_0_row_0(net156), .OUTPUT_1_row_0(net156));
	TSMC350nm_TA2Cell_Weak I__7 (.island_num(0), .row(7), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net232[0]), .VD_P_1_row_0(net233[0]), .VIN1_PLUSrow_0(net156), .VIN1_MINUSrow_0(net195), .VIN2_PLUSrow_0(net195), .VIN2_MINUSrow_0(net300), .OUTPUT_0_row_0(net195), .OUTPUT_1_row_0(net300));
	TSMC350nm_TA2Cell_Weak I__8 (.island_num(0), .row(8), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net234[0]), .VD_P_1_row_0(net235[0]), .VIN1_PLUSrow_0(net195), .VIN1_MINUSrow_0(net196), .VIN2_PLUSrow_0(net196), .VIN2_MINUSrow_0(net296), .OUTPUT_0_row_0(net196), .OUTPUT_1_row_0(net196));
	TSMC350nm_TA2Cell_Weak I__9 (.island_num(0), .row(9), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net236[0]), .VD_P_1_row_0(net237[0]), .VIN1_PLUSrow_0(net196), .VIN1_MINUSrow_0(net296), .VIN2_PLUSrow_0(net296), .VIN2_MINUSrow_0(net301), .OUTPUT_0_row_0(net296), .OUTPUT_1_row_0(net301), .VINJ_brow_0(net315), .GND_brow_0(net314));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5), .decode_n0_VINJ(net315), .decode_n0_GND(net314), .decode_n0_IN_0_(net308), .decode_n0_IN_1_(net309), .decode_n0_IN_2_(net310), .decode_n0_IN_3_(net311), .decode_n0_IN_4_(net312), .decode_n0_ENABLE(net313));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select), .switch_n0_prog_drainrail(net307), .switch_n0_VINJ(net315), .switch_n0_GND(net314));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch), .switch_n0_PR_0_(net218[0]), .switch_n0_PR_1_(net219[0]), .switch_n0_PR_2_(net220[0]), .switch_n0_PR_3_(net221[0]), .switch_n1_PR_0_(net222[0]), .switch_n1_PR_1_(net223[0]), .switch_n1_PR_2_(net224[0]), .switch_n1_PR_3_(net225[0]), .switch_n2_PR_0_(net226[0]), .switch_n2_PR_1_(net227[0]), .switch_n2_PR_2_(net228[0]), .switch_n2_PR_3_(net229[0]), .switch_n3_PR_0_(net230[0]), .switch_n3_PR_1_(net231[0]), .switch_n3_PR_2_(net232[0]), .switch_n3_PR_3_(net233[0]), .switch_n4_PR_0_(net234[0]), .switch_n4_PR_1_(net235[0]), .switch_n4_PR_2_(net236[0]), .switch_n4_PR_3_(net237[0]), .switch_n0_VDD(net315), .switch_n0_GND(net314), .switch_n0_RUN(net321));
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(2), .decode_n0_ENABLE(net304), .decode_n0_VINJV(net316), .decode_n0_GNDV(net317), .decode_n0_IN_0_(net305), .decode_n0_IN_1_(net306));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(1), .switch_n0_GND_T(net317), .switch_n0_VINJ_T(net316), .switch_n0_CTRL_B_0_(net293), .switch_n0_CTRL_B_1_(net294), .switch_n0_Vg_0_(net291), .switch_n0_Vg_1_(net292));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(0), .direction(horizontal), .col(0), .RUN_IN_0_(net302), .RUN_IN_1_(net302), .PROG(net320), .RUN(net321), .Vgsel(net303));


	/* Frame */ 
	tile_analog_frame cab_frame(.pin_layer(METAL3), .W_w_Vin(net295), .E_e_Vout(net296), .E_e_Vout_Buf_0_(net297), .E_e_Vout_Buf_1_(net298), .E_e_Vout_Buf_2_(net299), .E_e_Vout_Buf_3_(net300), .E_e_Vout_Buf_4_(net301), .N_n_Prog(net320), .N_n_Prog(net321), .N_n_VGRUN(net302), .N_n_VGPROG(net303), .N_n_VTUN(net318), .N_n_AVDD(net319), .N_n_gnd(net317), .S_s_gnd(net314), .N_n_vinj(net316), .S_s_vinj(net315), .S_s_Drainline_Prog(net307), .N_n_GateEnable(net304), .W_w_GateB_0_(net305), .W_w_GateB_1_(net306), .W_w_DrainEnable(net313), .W_w_DrainB_0_(net308), .W_w_DrainB_1_(net309), .W_w_DrainB_2_(net310), .W_w_DrainB_3_(net311), .W_w_DrainB_4_(net312));
 endmodule