VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER routingPitch REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.01 ;
LAYER POLY1
  TYPE MASTERSLICE ;
END POLY1

LAYER CONT
  TYPE CUT ;
  SPACING 0.4 ;
END CONT

LAYER METAL1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.5 ;
  SPACING 0.45 ;
  PROPERTY routingPitch 1.25 ;
END METAL1

LAYER VIA12
  TYPE CUT ;
  SPACING 0.45 ;
END VIA12

LAYER METAL2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.4 ;
END METAL2

LAYER VIA23
  TYPE CUT ;
  SPACING 0.45 ;
END VIA23

LAYER METAL3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.25 ;
END METAL3

LAYER VIA34
  TYPE CUT ;
  SPACING 0.45 ;
END VIA34

LAYER METAL4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.6 ;
  PROPERTY routingPitch 1.4 ;
END METAL4

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIARULE M4_M3 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL4 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1

VIARULE M1_POLY1 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 1 ;
END M1_POLY1

VIA M1_POLY1
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER POLY1 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.35 -0.35 0.35 0.35 ;
END M1_POLY1

VIA M2_M1
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL2 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M2_M1

VIA M3_M2
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL3 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL2 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M3_M2

VIA M4_M3
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL3 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M4_M3


MACRO TSMC350nm_4x2_Direct
  PIN Vd_l<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 20.3 0.7 20.8 ;
    END
  END Vd_l<0>
  PIN Vd_l<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 14.7 0.7 15.2 ;
    END
  END Vd_l<1>
  PIN Vd_l<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 7.0 0.7 7.5 ;
    END
  END Vd_l<2>
  PIN Vd_l<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 2.1 0.7 2.6 ;
    END
  END Vd_l<3>
  PIN Vd<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.2 2.1 21.0 2.6 ;
    END
  END Vd<3>
  PIN Vd<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.2 20.3 21.0 20.8 ;
    END
  END Vd<0>
  PIN Vd<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.2 7.0 21.0 7.5 ;
    END
  END Vd<2>
  PIN Vd<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.2 14.7 21.0 15.2 ;
    END
  END Vd<1>
  PIN GND<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 12.6 21.53 13.2 22.0 ;
    END
  END GND<1>
  PIN Vg<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 14.7 21.53 15.3 22.0 ;
    END
  END Vg<1>
  PIN VINJ<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 16.8 21.53 17.4 22.0 ;
    END
  END VINJ<1>
  PIN Vs<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 2.1 21.53 2.7 22.0 ;
    END
  END Vs<0>
  PIN Vg<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.3 21.53 6.9 22.0 ;
    END
  END Vg<0>
  PIN Vs<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 18.9 21.53 19.5 22.0 ;
    END
  END Vs<1>
  PIN VTUN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 10.5 21.53 11.1 22.0 ;
    END
  END VTUN
  PIN VINJ<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 4.2 21.53 4.8 22.0 ;
    END
  END VINJ<0>
  PIN GND<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 8.4 21.53 9.0 22.0 ;
    END
  END GND<0>
END TSMC350nm_4x2_Direct

END LIBRARY