module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(7), .GND_b_1_row_4(net2188[0:7]), .Vs_b_0_row_4(net124[0:7]), .Vs_b_1_row_4(net125[0:7]), .VINJ_b_1_row_4(net2195[0:7]), .Vsel_b_0_row_4(net2153[0:7]), .Vsel_b_1_row_4(net2154[0:7]), .Vg_b_0_row_4(net2167[0:7]), .Vg_b_1_row_4(net2168[0:7]), .VTUN_brow_4(net2181[0:7]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(17), .matrix_row(5), .matrix_col(9), .GND_b_1_row_4(net2231[0:9]), .Vs_b_0_row_4(net325[0:9]), .Vs_b_1_row_4(net326[0:9]), .VINJ_b_1_row_4(net2230[0:9]), .Vsel_b_0_row_4(net2232[0:9]), .Vsel_b_1_row_4(net2234[0:9]), .Vg_b_0_row_4(net2233[0:9]), .Vg_b_1_row_4(net2235[0:9]), .VTUN_brow_4(net2229[0:9]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(26), .matrix_row(5), .matrix_col(1), .A_0_col_0(net2569[0:5]), .A_1_col_0(net2570[0:5]), .A_2_col_0(net2571[0:5]), .A_3_col_0(net2572[0:5]), .Prog_brow_4(net2528[0:1]), .VDD_brow_4(net2507[0:1]), .GND_brow_4(net2231[8:9]), .Progrow_0(net2528[0:1]));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2208[0:1]), .Vsel_b_0_row_4(net2211[0:1]), .Vsel_b_1_row_4(net2212[0:1]), .Vg_b_0_row_4(net2213[0:1]), .Vg_b_1_row_4(net2214[0:1]), .VTUN_brow_4(net2209[0:1]), .GND_b_1_row_4(net2210[0:1]));
	S_BLOCK_BUFFER I__4 (.island_num(0), .row(0), .col(8), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__5 (.island_num(0), .row(0), .col(9), .matrix_row(4), .matrix_col(1), .n_0_row_0(net2476[0:1]), .n_1_row_0(net2477[0:1]), .n_2_row_0(net2478[0:1]), .n_3_row_0(net2479[0:1]));
	S_BLOCK_CONN_PINS I__6 (.island_num(0), .row(4), .col(9), .matrix_row(1), .matrix_col(1), .s_0_row_0(net2508), .s_1_row_0(net2509), .s_2_row_0(net2510), .s_3_row_0(net2511));
	S_BLOCK_SPACE_UP_PINS I__7 (.island_num(0), .row(0), .col(10), .matrix_row(3), .matrix_col(1), .n_0_row_0(net2480[0:1]), .n_1_row_0(net2481[0:1]), .n_2_row_0(net2482[0:1]), .n_3_row_0(net2483[0:1]));
	S_BLOCK_CONN_PINS I__8 (.island_num(0), .row(3), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__9 (.island_num(0), .row(4), .col(10), .matrix_row(1), .matrix_col(1), .s_0_row_0(net2512), .s_1_row_0(net2513), .s_2_row_0(net2514), .s_3_row_0(net2515));
	S_BLOCK_SPACE_UP_PINS I__10 (.island_num(0), .row(0), .col(11), .matrix_row(2), .matrix_col(1), .n_0_row_0(net2484[0:1]), .n_1_row_0(net2485[0:1]), .n_2_row_0(net2486[0:1]), .n_3_row_0(net2487[0:1]));
	S_BLOCK_CONN_PINS I__11 (.island_num(0), .row(2), .col(11), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__12 (.island_num(0), .row(3), .col(11), .matrix_row(2), .matrix_col(1), .s_0_row_1(net2516[0:1]), .s_1_row_1(net2517[0:1]), .s_2_row_1(net2518[0:1]), .s_3_row_1(net2519[0:1]));
	S_BLOCK_SPACE_UP_PINS I__13 (.island_num(0), .row(0), .col(12), .matrix_row(1), .matrix_col(1), .n_0_row_0(net2488), .n_1_row_0(net2489), .n_2_row_0(net2490), .n_3_row_0(net2491));
	S_BLOCK_CONN_PINS I__14 (.island_num(0), .row(1), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__15 (.island_num(0), .row(2), .col(12), .matrix_row(3), .matrix_col(1), .s_0_row_2(net2520[0:1]), .s_1_row_2(net2521[0:1]), .s_2_row_2(net2522[0:1]), .s_3_row_2(net2523[0:1]));
	S_BLOCK_CONN_PINS I__16 (.island_num(0), .row(0), .col(13), .matrix_row(1), .matrix_col(1), .n_0_row_0(net2492), .n_1_row_0(net2493), .n_2_row_0(net2494), .n_3_row_0(net2495));
	S_BLOCK_SPACE_DOWN_PINS I__17 (.island_num(0), .row(1), .col(13), .matrix_row(4), .matrix_col(1), .s_0_row_3(net2524[0:1]), .s_1_row_3(net2525[0:1]), .s_2_row_3(net2526[0:1]), .s_3_row_3(net2527[0:1]));
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2215[0:1]), .Vsel_b_0_row_4(net2218[0:1]), .Vsel_b_1_row_4(net2219[0:1]), .Vg_b_0_row_4(net2220[0:1]), .Vg_b_1_row_4(net2221[0:1]), .VTUN_brow_4(net2216[0:1]), .GND_b_1_row_4(net2217[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2222[0:1]), .Vsel_b_0_row_4(net2225[0:1]), .Vsel_b_1_row_4(net2226[0:1]), .Vg_b_0_row_4(net2227[0:1]), .Vg_b_1_row_4(net2228[0:1]), .VTUN_brow_4(net2223[0:1]), .GND_b_1_row_4(net2224[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(6), .decode_n2_VGRUN_0_(net2472[0]), .decode_n2_VGRUN_1_(net2473[0]), .decode_n2_VGRUN_2_(net2474[0]), .decode_n2_VGRUN_3_(net2475[0]), .decode_n7_VGRUN_2_(net2555[0]), .decode_n7_VGRUN_3_(net2556[0]), .decode_n8_VGRUN_0_(net2557[0]), .decode_n8_VGRUN_1_(net2558[0]), .decode_n4_n0_RUN_OUT_0_(net2302), .decode_n4_n0_RUN_OUT_1_(net2303), .decode_n4_n0_RUN_OUT_2_(net2308), .decode_n4_n0_RUN_OUT_3_(net2309), .decode_n4_n1_RUN_OUT_0_(net2314), .decode_n4_n1_RUN_OUT_1_(net2315), .decode_n4_n1_RUN_OUT_2_(net2320), .decode_n4_n1_RUN_OUT_3_(net2321), .decode_n4_n2_RUN_OUT_0_(net2326), .decode_n4_n2_RUN_OUT_1_(net2327), .decode_n4_n2_RUN_OUT_2_(net2332), .decode_n4_n2_RUN_OUT_3_(net2333), .decode_n4_n3_RUN_OUT_0_(net2338), .decode_n4_n3_RUN_OUT_1_(net2339), .decode_n4_n3_RUN_OUT_2_(net2344), .decode_n4_n3_RUN_OUT_3_(net2345), .decode_n4_n0_OUT_0_(net2300), .decode_n4_n0_OUT_1_(net2301), .decode_n4_n0_OUT_2_(net2306), .decode_n4_n0_OUT_3_(net2307), .decode_n4_n1_OUT_0_(net2312), .decode_n4_n1_OUT_1_(net2313), .decode_n4_n1_OUT_2_(net2318), .decode_n4_n1_OUT_3_(net2319), .decode_n4_n2_OUT_0_(net2324), .decode_n4_n2_OUT_1_(net2325), .decode_n4_n2_OUT_2_(net2330), .decode_n4_n2_OUT_3_(net2331), .decode_n4_n3_OUT_0_(net2336), .decode_n4_n3_OUT_1_(net2337), .decode_n4_n3_OUT_2_(net2342), .decode_n4_n3_OUT_3_(net2343), .decode_n4_n4_OUT_0_(net2348), .decode_n4_n4_OUT_1_(net2349), .decode_n4_n5_OUT_0_(net2352), .decode_n4_n5_OUT_1_(net2353), .decode_n4_n5_OUT_2_(net2356), .decode_n4_n5_OUT_3_(net2357), .decode_n4_n6_OUT_0_(net2360), .decode_n4_n6_OUT_1_(net2361), .decode_n4_n6_OUT_2_(net2364), .decode_n4_n6_OUT_3_(net2365), .decode_n4_n7_OUT_0_(net2368), .decode_n4_n7_OUT_1_(net2369), .decode_n4_n7_OUT_2_(net2372), .decode_n4_n7_OUT_3_(net2373), .decode_n4_n8_OUT_0_(net2376), .decode_n4_n8_OUT_1_(net2377), .decode_n4_n8_OUT_2_(net2380), .decode_n4_n8_OUT_3_(net2381), .decode_n4_n9_OUT_0_(net2384), .decode_n4_n9_OUT_1_(net2385), .decode_n4_n9_OUT_2_(net2388), .decode_n4_n9_OUT_3_(net2389), .decode_n0_ENABLE(net2496), .decode_n4_n0_VINJ_b_0_(net2298), .decode_n4_n0_VINJ_b_1_(net2304), .decode_n4_n1_VINJ_b_0_(net2310), .decode_n4_n1_VINJ_b_1_(net2316), .decode_n4_n2_VINJ_b_0_(net2322), .decode_n4_n2_VINJ_b_1_(net2328), .decode_n4_n3_VINJ_b_0_(net2334), .decode_n4_n3_VINJ_b_1_(net2340), .decode_n4_n4_VINJ_b_0_(net2346), .decode_n4_n5_VINJ_b_0_(net2350), .decode_n4_n5_VINJ_b_1_(net2354), .decode_n4_n6_VINJ_b_0_(net2358), .decode_n4_n6_VINJ_b_1_(net2362), .decode_n4_n7_VINJ_b_0_(net2366), .decode_n4_n7_VINJ_b_1_(net2370), .decode_n4_n8_VINJ_b_0_(net2374), .decode_n4_n8_VINJ_b_1_(net2378), .decode_n4_n9_VINJ_b_0_(net2382), .decode_n4_n9_VINJ_b_1_(net2386), .decode_n4_n0_GND_b_0_(net2299), .decode_n4_n0_GND_b_1_(net2305), .decode_n4_n1_GND_b_0_(net2311), .decode_n4_n1_GND_b_1_(net2317), .decode_n4_n2_GND_b_0_(net2323), .decode_n4_n2_GND_b_1_(net2329), .decode_n4_n3_GND_b_0_(net2335), .decode_n4_n3_GND_b_1_(net2341), .decode_n4_n4_GND_b_0_(net2347), .decode_n4_n5_GND_b_0_(net2351), .decode_n4_n5_GND_b_1_(net2355), .decode_n4_n6_GND_b_0_(net2359), .decode_n4_n6_GND_b_1_(net2363), .decode_n4_n7_GND_b_0_(net2367), .decode_n4_n7_GND_b_1_(net2371), .decode_n4_n8_GND_b_0_(net2375), .decode_n4_n8_GND_b_1_(net2379), .decode_n4_n9_GND_b_0_(net2383), .decode_n4_n9_GND_b_1_(net2387), .decode_n0_VINJV(net2503), .decode_n0_GNDV(net2505));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(26), .switch_n0_VPWR_0_(net2302), .switch_n0_VPWR_1_(net2303), .switch_n1_VPWR_0_(net2308), .switch_n1_VPWR_1_(net2309), .switch_n2_VPWR_0_(net2314), .switch_n2_VPWR_1_(net2315), .switch_n3_VPWR_0_(net2320), .switch_n3_VPWR_1_(net2321), .switch_n4_VPWR_0_(net2326), .switch_n4_VPWR_1_(net2327), .switch_n5_VPWR_0_(net2332), .switch_n5_VPWR_1_(net2333), .switch_n6_VPWR_0_(net2338), .switch_n6_VPWR_1_(net2339), .switch_n7_VPWR_0_(net2344), .switch_n7_VPWR_1_(net2345), .switch_n0_RUN_IN_0_(net2559[0]), .switch_n0_RUN_IN_1_(net2559[0]), .switch_n1_RUN_IN_0_(net2559[0]), .switch_n1_RUN_IN_1_(net2559[0]), .switch_n2_RUN_IN_0_(net2559[0]), .switch_n2_RUN_IN_1_(net2559[0]), .switch_n3_RUN_IN_0_(net2559[0]), .switch_n3_RUN_IN_1_(net2559[0]), .switch_n4_RUN_IN_0_(net2559[0]), .switch_n4_RUN_IN_1_(net2559[0]), .switch_n5_RUN_IN_0_(net2559[0]), .switch_n5_RUN_IN_1_(net2559[0]), .switch_n6_RUN_IN_0_(net2559[0]), .switch_n6_RUN_IN_1_(net2559[0]), .switch_n7_RUN_IN_0_(net2559[0]), .switch_n7_RUN_IN_1_(net2559[0]), .switch_n14_RUN_IN_0_(net2559[0]), .switch_n14_RUN_IN_1_(net2559[0]), .switch_n16_RUN_IN_0_(net2559[0]), .switch_n16_RUN_IN_1_(net2559[0]), .switch_n17_RUN_IN_0_(net2559[0]), .switch_n17_RUN_IN_1_(net2559[0]), .switch_n18_RUN_IN_0_(net2559[0]), .switch_n18_RUN_IN_1_(net2559[0]), .switch_n19_RUN_IN_0_(net2559[0]), .switch_n19_RUN_IN_1_(net2559[0]), .switch_n20_RUN_IN_0_(net2559[0]), .switch_n20_RUN_IN_1_(net2559[0]), .switch_n21_RUN_IN_0_(net2559[0]), .switch_n21_RUN_IN_1_(net2559[0]), .switch_n22_RUN_IN_0_(net2559[0]), .switch_n22_RUN_IN_1_(net2559[0]), .switch_n23_RUN_IN_0_(net2559[0]), .switch_n23_RUN_IN_1_(net2559[0]), .switch_n24_RUN_IN_0_(net2559[0]), .switch_n24_RUN_IN_1_(net2559[0]), .switch_n25_RUN_IN_0_(net2559[0]), .switch_n25_RUN_IN_1_(net2559[0]), .switch_n0_GND_T(net2299), .switch_n1_GND_T(net2305), .switch_n2_GND_T(net2311), .switch_n3_GND_T(net2317), .switch_n4_GND_T(net2323), .switch_n5_GND_T(net2329), .switch_n6_GND_T(net2335), .switch_n7_GND_T(net2341), .switch_n14_GND_T(net2347), .switch_n16_GND_T(net2351), .switch_n17_GND_T(net2355), .switch_n18_GND_T(net2359), .switch_n19_GND_T(net2363), .switch_n20_GND_T(net2367), .switch_n21_GND_T(net2371), .switch_n22_GND_T(net2375), .switch_n23_GND_T(net2379), .switch_n24_GND_T(net2383), .switch_n25_GND_T(net2387), .switch_n0_VTUN_T(net2560[0]), .switch_n0_decode_0_(net2300), .switch_n0_decode_1_(net2301), .switch_n1_decode_0_(net2306), .switch_n1_decode_1_(net2307), .switch_n2_decode_0_(net2312), .switch_n2_decode_1_(net2313), .switch_n3_decode_0_(net2318), .switch_n3_decode_1_(net2319), .switch_n4_decode_0_(net2324), .switch_n4_decode_1_(net2325), .switch_n5_decode_0_(net2330), .switch_n5_decode_1_(net2331), .switch_n6_decode_0_(net2336), .switch_n6_decode_1_(net2337), .switch_n7_decode_0_(net2342), .switch_n7_decode_1_(net2343), .switch_n14_decode_0_(net2348), .switch_n14_decode_1_(net2349), .switch_n16_decode_0_(net2352), .switch_n16_decode_1_(net2353), .switch_n17_decode_0_(net2356), .switch_n17_decode_1_(net2357), .switch_n18_decode_0_(net2360), .switch_n18_decode_1_(net2361), .switch_n19_decode_0_(net2364), .switch_n19_decode_1_(net2365), .switch_n20_decode_0_(net2368), .switch_n20_decode_1_(net2369), .switch_n21_decode_0_(net2372), .switch_n21_decode_1_(net2373), .switch_n22_decode_0_(net2376), .switch_n22_decode_1_(net2377), .switch_n23_decode_0_(net2380), .switch_n23_decode_1_(net2381), .switch_n24_decode_0_(net2384), .switch_n24_decode_1_(net2385), .switch_n25_decode_0_(net2388), .switch_n25_decode_1_(net2389), .switch_n0_VINJ_T(net2298), .switch_n1_VINJ_T(net2304), .switch_n2_VINJ_T(net2310), .switch_n3_VINJ_T(net2316), .switch_n4_VINJ_T(net2322), .switch_n5_VINJ_T(net2328), .switch_n6_VINJ_T(net2334), .switch_n7_VINJ_T(net2340), .switch_n14_VINJ_T(net2346), .switch_n16_VINJ_T(net2350), .switch_n17_VINJ_T(net2354), .switch_n18_VINJ_T(net2358), .switch_n19_VINJ_T(net2362), .switch_n20_VINJ_T(net2366), .switch_n21_VINJ_T(net2370), .switch_n22_VINJ_T(net2374), .switch_n23_VINJ_T(net2378), .switch_n24_VINJ_T(net2382), .switch_n25_VINJ_T(net2386), .switch_n0_RUN(net2529), .switch_n0_vgsel_r(net2530));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5), .decode_n0_IN_0_(net2568), .decode_n0_IN_1_(net2567), .decode_n0_IN_2_(net2566), .decode_n0_IN_3_(net2565), .decode_n0_IN_4_(net2564), .decode_n0_ENABLE(net2595));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select), .switch_n0_prog_drainrail(net2497), .switch_n0_run_drainrail(net2498), .switch_n0_VINJ(net2504), .switch_n0_GND(net2506));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch), .switch_n0_In_0_(net2535[0]), .switch_n0_In_1_(net2536[0]), .switch_n0_In_2_(net2537[0]), .switch_n0_In_3_(net2538[0]), .switch_n1_In_0_(net2539[0]), .switch_n1_In_1_(net2540[0]), .switch_n1_In_2_(net2541[0]), .switch_n1_In_3_(net2542[0]), .switch_n2_In_0_(net2543[0]), .switch_n2_In_1_(net2544[0]), .switch_n2_In_2_(net2545[0]), .switch_n2_In_3_(net2546[0]), .switch_n3_In_0_(net2547[0]), .switch_n3_In_1_(net2548[0]), .switch_n3_In_2_(net2549[0]), .switch_n3_In_3_(net2550[0]), .switch_n4_In_0_(net2551[0]), .switch_n4_In_1_(net2552[0]), .switch_n4_In_2_(net2553[0]), .switch_n4_In_3_(net2554[0]), .switch_n0_VDD(net2504), .switch_n0_GND(net2506), .switch_n0_RUN(net2529));
	none switch_ind(.island_num(0), .direction(horizontal), .col(8));
	none switch_ind(.island_num(0), .direction(horizontal), .col(9));
	none switch_ind(.island_num(0), .direction(horizontal), .col(10));
	none switch_ind(.island_num(0), .direction(horizontal), .col(11));
	none switch_ind(.island_num(0), .direction(horizontal), .col(12));
	none switch_ind(.island_num(0), .direction(horizontal), .col(13));
	none switch_ind(.island_num(0), .direction(horizontal), .col(15));


	/* Island 1 */
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__0 (.island_num(1), .row(0), .col(0), .matrix_row(1), .matrix_col(8));
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(7), .matrix_col(8), .GND_b_0_row_6(net1181[0:8]), .GND_b_1_row_6(net1182[0:8]), .Vs_b_0_row_6(net1191[0:8]), .Vs_b_1_row_6(net1192[0:8]), .VINJ_b_0_row_6(net1195[0:8]), .VINJ_b_1_row_6(net1196[0:8]), .Vsel_b_0_row_6(net1199[0:8]), .Vsel_b_1_row_6(net1200[0:8]), .Vg_b_0_row_6(net1203[0:8]), .Vg_b_1_row_6(net1204[0:8]), .VTUN_brow_6(net1207[0:8]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(8), .matrix_row(6), .matrix_col(10));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(7), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2055), .P_1_row_0(net2056), .A_0_row_0(net2057), .A_1_row_0(net2058), .A_2_row_0(net2059), .A_3_row_0(net2060));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2067), .P_1_row_0(net2068), .A_0_row_0(net2069), .A_1_row_0(net2070), .A_2_row_0(net2071), .A_3_row_0(net2072));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2085), .P_1_row_0(net2086), .A_0_row_0(net2087), .A_1_row_0(net2088), .A_2_row_0(net2089), .A_3_row_0(net2090));
	TSMC350nm_4TGate_ST_BMatrix_NoSwitch I__8 (.island_num(1), .row(3), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2103), .P_1_row_0(net2104), .P_2_row_0(net2105), .P_3_row_0(net2106), .A_0_row_0(net2107), .A_1_row_0(net2108), .A_2_row_0(net2109), .A_3_row_0(net2110));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2122), .P_1_row_0(net2123), .P_2_row_0(net2124), .P_3_row_0(net2125), .A_0_row_0(net2126), .A_1_row_0(net2127));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net2137), .A_1_row_0(net2138), .A_2_row_0(net2139), .A_3_row_0(net2140));
	TSMC350nm_4TGate_ST_BMatrix I__11 (.island_num(1), .row(6), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net2144), .A_1_row_0(net2145), .A_2_row_0(net2146), .A_3_row_0(net2147));
	TSMC350nm_4TGate_ST_BMatrix I__12 (.island_num(1), .row(7), .col(18), .matrix_row(1), .matrix_col(1), .Prog_brow_0(net2471[0]), .VDD_brow_0(net2507[0]), .GND_brow_0(net2231[8]));
	TSMC350nm_OutMtrx_IndrctSwcs I__13 (.island_num(1), .row(9), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__14 (.island_num(1), .row(10), .col(8), .matrix_row(2), .matrix_col(10), .Vd_Rl_0_col_0(net1902[0:2]), .Vd_Rl_1_col_0(net1903[0:2]), .Vd_Rl_2_col_0(net1904[0:2]), .Vd_Rl_3_col_0(net1905[0:2]), .Vd_Pl_0_col_0(net1906[0:2]), .Vd_Pl_1_col_0(net1907[0:2]), .Vd_Pl_2_col_0(net1908[0:2]), .Vd_Pl_3_col_0(net1909[0:2]));
	TSMC350nm_4TGate_ST_BMatrix I__15 (.island_num(1), .row(10), .col(18), .matrix_row(2), .matrix_col(1), .A_0_col_0(net2499[0:2]), .A_1_col_0(net2500[0:2]), .A_2_col_0(net2501[0:2]), .A_3_col_0(net2502[0:2]), .Prog_brow_1(net2471[0:1]), .VDD_brow_1(net2507[0:1]), .GND_brow_1(net2231[8:9]));
	TSMC350nm_TA2Cell_Weak cab_device_16 (.island_num(1), .row(2), .col(19), .VD_P_0_(net2055), .VD_P_1_(net2056), .VIN1_PLUS(net2057), .VIN1_MINUS(net2058), .VIN2_PLUS(net2059), .VIN2_MINUS(net2060), .OUTPUT_0_(net2061[0]), .OUTPUT_1_(net2062[0]), .Vsel_0_(net2131), .Vsel_1_(net2132), .RUN(net2063), .Vg_0_(net2133), .Vg_1_(net2134), .PROG(net2528[0]), .VTUN(net2064), .VINJ(net2065), .GND(net2066), .VPWR(net2563[0]), .Vsel_b_0_(net2075), .Vsel_b_1_(net2076), .RUN_b(net2077), .Vg_b_0_(net2078), .Vg_b_1_(net2079), .PROG_b(net2080), .VTUN_b(net2081), .VINJ_b(net2082), .GND_b(net2083), .VPWR_b(net2084));
	TSMC350nm_TA2Cell_Weak cab_device_17 (.island_num(1), .row(3), .col(19), .VD_P_0_(net2067), .VD_P_1_(net2068), .VIN1_PLUS(net2069), .VIN1_MINUS(net2070), .VIN2_PLUS(net2071), .VIN2_MINUS(net2072), .OUTPUT_0_(net2073[0]), .OUTPUT_1_(net2074[0]), .Vsel_0_(net2075), .Vsel_1_(net2076), .RUN(net2077), .Vg_0_(net2078), .Vg_1_(net2079), .PROG(net2080), .VTUN(net2081), .VINJ(net2082), .GND(net2083), .VPWR(net2084), .Vsel_b_0_(net2093), .Vsel_b_1_(net2094), .RUN_b(net2095), .Vg_b_0_(net2096), .Vg_b_1_(net2097), .PROG_b(net2098), .VTUN_b(net2099), .VINJ_b(net2100), .GND_b(net2101), .VPWR_b(net2102));
	TSMC350nm_TA2Cell_Strong cab_device_18 (.island_num(1), .row(4), .col(19), .VD_P_0_(net2085), .VD_P_1_(net2086), .VIN1_PLUS(net2087), .VIN1_MINUS(net2088), .VIN2_PLUS(net2089), .VIN2_MINUS(net2090), .OUTPUT_0_(net2091[0]), .OUTPUT_1_(net2092[0]), .Vsel_0_(net2093), .Vsel_1_(net2094), .RUN(net2095), .Vg_0_(net2096), .Vg_1_(net2097), .PROG(net2098), .VTUN(net2099), .VINJ(net2100), .GND(net2101), .VPWR(net2102), .Vg_b_0_(net2118), .PROG_b(net2121), .VTUN_b(net2119), .VINJ_b(net2117), .GND_b(net2120));
	TSMC350nm_4WTA_IndirectProg cab_device_19 (.island_num(1), .row(5), .col(19), .VD_P_0_(net2103), .VD_P_1_(net2104), .VD_P_2_(net2105), .VD_P_3_(net2106), .Iin_0_(net2107), .Iin_1_(net2108), .Iin_2_(net2109), .Iin_3_(net2110), .Vout_0_(net2111[0]), .Vout_1_(net2112[0]), .Vout_2_(net2113[0]), .Vout_3_(net2114[0]), .Vmid(net2115[0]), .Vbias(net2116[0]), .Vsel(net2131), .Vs(net2563[0]), .VINJ(net2117), .Vg(net2118), .VTUN(net2119), .GND(net2120), .PROG(net2121), .VINJ_b(net2130), .VTUN_b(net2136), .GND_b(net2135));
	TSMC350nm_Cap_Bank cab_device_20 (.island_num(1), .row(6), .col(19), .VD_P_0_(net2122), .VD_P_1_(net2123), .VD_P_2_(net2124), .VD_P_3_(net2125), .VIN_0_(net2126), .VIN_1_(net2127), .OUT_0_(net2128[0]), .OUT_1_(net2129[0]), .VINJ(net2130), .Vsel_0_(net2131), .Vsel_1_(net2132), .Vg_0_(net2133), .Vg_1_(net2134), .GND(net2135), .VTUN(net2136), .GND_b(net2143));
	TSMC350nm_NandPfets cab_device_21 (.island_num(1), .row(7), .col(19), .GATE_N(net2137), .SOURCE_N(net2138), .GATE_P(net2139), .SOURCE_P(net2140), .DRAIN_N(net2141[0]), .DRAIN_P(net2142[0]), .VPWR(net2563[0]), .GND(net2143), .VPWR_b(net2151), .GND_b(net2152));
	TSMC350nm_TGate_2nMirror cab_device_22 (.island_num(1), .row(8), .col(19), .IN_CM_0_(net2144), .IN_CM_1_(net2145), .SelN(net2146), .IN_TG(net2147), .OUT_CM_0_(net2148[0]), .OUT_CM_1_(net2149[0]), .OUT_TG(net2150[0]), .VPWR(net2151), .GND(net2152));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6), .decode_n0_IN_0_(net2594), .decode_n0_IN_1_(net2593), .decode_n0_IN_2_(net2592), .decode_n0_IN_3_(net2591), .decode_n0_IN_4_(net2590), .decode_n0_IN_5_(net2589), .decode_n0_ENABLE(net2595));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(1), .direction(vertical), .num(12), .type(drain_select), .switch_n0_prog_drainrail(net2497), .switch_n0_run_drainrail(net2498));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(12), .type(prog_switch), .switch_n8_PR_0_(net2455[0]), .switch_n8_PR_1_(net2459[0]), .switch_n8_PR_2_(net2463[0]), .switch_n8_PR_3_(net2467[0]), .switch_n8_In_0_(net2454[0]), .switch_n8_In_1_(net2458[0]), .switch_n8_In_2_(net2462[0]), .switch_n8_In_3_(net2466[0]), .switch_n0_RUN(net2529));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(20), .switch_n0_Input_0_(net2507[0]), .switch_n0_Input_1_(net2188[0]), .switch_n1_Input_0_(net124[1]), .switch_n1_Input_1_(net125[1]), .switch_n2_Input_0_(net124[2]), .switch_n2_Input_1_(net125[2]), .switch_n3_Input_0_(net124[3]), .switch_n3_Input_1_(net125[3]), .switch_n4_Input_0_(net325[0]), .switch_n4_Input_1_(net326[0]), .switch_n5_Input_0_(net325[1]), .switch_n5_Input_1_(net326[1]), .switch_n6_Input_0_(net325[2]), .switch_n6_Input_1_(net326[2]), .switch_n7_Input_0_(net325[3]), .switch_n7_Input_1_(net326[3]), .switch_n8_Input_0_(net2453[0]), .switch_n8_Input_1_(net2061[0]), .switch_n9_Input_0_(net2062[0]), .switch_n9_Input_1_(net2073[0]), .switch_n10_Input_0_(net2074[0]), .switch_n10_Input_1_(net2091[0]), .switch_n11_Input_0_(net2092[0]), .switch_n11_Input_1_(net2111[0]), .switch_n12_Input_0_(net2112[0]), .switch_n12_Input_1_(net2113[0]), .switch_n13_Input_0_(net2114[0]), .switch_n13_Input_1_(net2115[0]), .switch_n14_Input_0_(net2116[0]), .switch_n14_Input_1_(net2128[0]), .switch_n15_Input_0_(net2129[0]), .switch_n15_Input_1_(net2141[0]), .switch_n16_Input_0_(net2142[0]), .switch_n16_Input_1_(net2148[0]), .switch_n17_Input_0_(net2149[0]), .switch_n17_Input_1_(net2150[0]), .switch_n0_GND(net2188[0]), .switch_n1_GND(net2188[1]), .switch_n2_GND(net2188[2]), .switch_n3_GND(net2188[3]), .switch_n4_GND(net2188[4]), .switch_n5_GND(net2188[5]), .switch_n6_GND(net2188[6]), .switch_n7_GND(net2210[0]), .switch_n8_GND(net2217[0]), .switch_n9_GND(net2224[0]), .switch_n10_GND(net2231[0]), .switch_n11_GND(net2231[1]), .switch_n12_GND(net2231[2]), .switch_n13_GND(net2231[3]), .switch_n14_GND(net2231[4]), .switch_n15_GND(net2231[5]), .switch_n16_GND(net2231[6]), .switch_n17_GND(net2231[7]), .switch_n18_GND(net2231[8]), .switch_n0_Vsel_0_(net2153[0]), .switch_n0_Vsel_1_(net2154[0]), .switch_n1_Vsel_0_(net2153[1]), .switch_n1_Vsel_1_(net2154[1]), .switch_n2_Vsel_0_(net2153[2]), .switch_n2_Vsel_1_(net2154[2]), .switch_n3_Vsel_0_(net2153[3]), .switch_n3_Vsel_1_(net2154[3]), .switch_n4_Vsel_0_(net2153[4]), .switch_n4_Vsel_1_(net2154[4]), .switch_n5_Vsel_0_(net2153[5]), .switch_n5_Vsel_1_(net2154[5]), .switch_n6_Vsel_0_(net2153[6]), .switch_n6_Vsel_1_(net2154[6]), .switch_n7_Vsel_0_(net2212[0]), .switch_n7_Vsel_1_(net2211[0]), .switch_n8_Vsel_0_(net2219[0]), .switch_n8_Vsel_1_(net2218[0]), .switch_n9_Vsel_0_(net2226[0]), .switch_n9_Vsel_1_(net2225[0]), .switch_n10_Vsel_0_(net2232[0]), .switch_n10_Vsel_1_(net2234[0]), .switch_n11_Vsel_0_(net2232[1]), .switch_n11_Vsel_1_(net2234[1]), .switch_n12_Vsel_0_(net2232[2]), .switch_n12_Vsel_1_(net2234[2]), .switch_n13_Vsel_0_(net2232[3]), .switch_n13_Vsel_1_(net2234[3]), .switch_n14_Vsel_0_(net2232[4]), .switch_n14_Vsel_1_(net2234[4]), .switch_n15_Vsel_0_(net2232[5]), .switch_n15_Vsel_1_(net2234[5]), .switch_n16_Vsel_0_(net2232[6]), .switch_n16_Vsel_1_(net2234[6]), .switch_n17_Vsel_0_(net2232[7]), .switch_n17_Vsel_1_(net2234[7]), .switch_n18_Vsel_0_(net2232[8]), .switch_n18_Vsel_1_(net2234[8]), .switch_n0_Vg_global_0_(net2167[0]), .switch_n0_Vg_global_1_(net2168[0]), .switch_n1_Vg_global_0_(net2167[1]), .switch_n1_Vg_global_1_(net2168[1]), .switch_n2_Vg_global_0_(net2167[2]), .switch_n2_Vg_global_1_(net2168[2]), .switch_n3_Vg_global_0_(net2167[3]), .switch_n3_Vg_global_1_(net2168[3]), .switch_n4_Vg_global_0_(net2167[4]), .switch_n4_Vg_global_1_(net2168[4]), .switch_n5_Vg_global_0_(net2167[5]), .switch_n5_Vg_global_1_(net2168[5]), .switch_n6_Vg_global_0_(net2167[6]), .switch_n6_Vg_global_1_(net2168[6]), .switch_n7_Vg_global_0_(net2214[0]), .switch_n7_Vg_global_1_(net2213[0]), .switch_n8_Vg_global_0_(net2221[0]), .switch_n8_Vg_global_1_(net2220[0]), .switch_n9_Vg_global_0_(net2228[0]), .switch_n9_Vg_global_1_(net2227[0]), .switch_n10_Vg_global_0_(net2233[0]), .switch_n10_Vg_global_1_(net2235[0]), .switch_n11_Vg_global_0_(net2233[1]), .switch_n11_Vg_global_1_(net2235[1]), .switch_n12_Vg_global_0_(net2233[2]), .switch_n12_Vg_global_1_(net2235[2]), .switch_n13_Vg_global_0_(net2233[3]), .switch_n13_Vg_global_1_(net2235[3]), .switch_n14_Vg_global_0_(net2233[4]), .switch_n14_Vg_global_1_(net2235[4]), .switch_n15_Vg_global_0_(net2233[5]), .switch_n15_Vg_global_1_(net2235[5]), .switch_n16_Vg_global_0_(net2233[6]), .switch_n16_Vg_global_1_(net2235[6]), .switch_n17_Vg_global_0_(net2233[7]), .switch_n17_Vg_global_1_(net2235[7]), .switch_n18_Vg_global_0_(net2233[8]), .switch_n18_Vg_global_1_(net2235[8]), .switch_n0_VTUN(net2181[0]), .switch_n1_VTUN(net2181[1]), .switch_n2_VTUN(net2181[2]), .switch_n3_VTUN(net2181[3]), .switch_n4_VTUN(net2181[4]), .switch_n5_VTUN(net2181[5]), .switch_n6_VTUN(net2181[6]), .switch_n7_VTUN(net2209[0]), .switch_n8_VTUN(net2216[0]), .switch_n9_VTUN(net2223[0]), .switch_n10_VTUN(net2229[0]), .switch_n11_VTUN(net2229[1]), .switch_n12_VTUN(net2229[2]), .switch_n13_VTUN(net2229[3]), .switch_n14_VTUN(net2229[4]), .switch_n15_VTUN(net2229[5]), .switch_n16_VTUN(net2229[6]), .switch_n17_VTUN(net2229[7]), .switch_n18_VTUN(net2229[8]), .switch_n0_VINJ(net2195[0]), .switch_n1_VINJ(net2195[1]), .switch_n2_VINJ(net2195[2]), .switch_n3_VINJ(net2195[3]), .switch_n4_VINJ(net2195[4]), .switch_n5_VINJ(net2195[5]), .switch_n6_VINJ(net2195[6]), .switch_n7_VINJ(net2208[0]), .switch_n8_VINJ(net2215[0]), .switch_n9_VINJ(net2222[0]), .switch_n10_VINJ(net2230[0]), .switch_n11_VINJ(net2230[1]), .switch_n12_VINJ(net2230[2]), .switch_n13_VINJ(net2230[3]), .switch_n14_VINJ(net2230[4]), .switch_n15_VINJ(net2230[5]), .switch_n16_VINJ(net2230[6]), .switch_n17_VINJ(net2230[7]), .switch_n18_VINJ(net2230[8]), .switch_n0_Vgrun_r(net2559[0]), .switch_n0_AVDD_r(net2563[0]), .switch_n0_run_r(net2470), .switch_n0_prog_r(net2471[0]), .switch_n0_run(net2529));
	none switch_ind(.island_num(1), .direction(horizontal), .col(18));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(19), .VPWR_0_(net2507[0]), .VPWR_1_(net2507[0]), .RUN_IN_0_(net2559[0]), .RUN_IN_1_(net2559[0]), .GND_T(net2231[8]), .VTUN_T(net2229[8]), .decode_0_(net2232[8]), .decode_1_(net2234[8]), .VINJ_T(net2230[8]), .GND(net2066), .CTRL_B_0_(net2131), .CTRL_B_1_(net2132), .run_r(net2063), .prog_r(net2528[0]), .Vg_0_(net2133), .Vg_1_(net2134), .VTUN(net2064), .VINJ(net2065), .VDD_1_(net2563[0]), .PROG(net2471[0]), .RUN(net2470), .Vgsel(net2530));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net1191[0:6]), .out_1_row_0(net1192[0:6]), .VINJ_0_row_0(net1195[0:6]), .VINJ_1_row_0(net1196[0:6]), .Vsel_0_row_0(net1199[0:6]), .Vsel_1_row_0(net1200[0:6]), .Vg_0_row_0(net1203[0:6]), .Vg_1_row_0(net1204[0:6]), .GNDrow_0(net1181[0:6]), .VTUNrow_0(net1207[0:6]), .Dcol_0(net124[6:7]), .CLKcol_0(net125[6:7]), .Qcol_5(net326[6:7]), .comcol_0(net2453[0:1]), .VDDcol_0(net2563[0:1]), .Vd_Pcol_0(net2467[0:1]), .Vd_in_0_col_0(net2454[0:1]), .Vd_in_1_col_0(net2458[0:1]), .Vd_in_2_col_0(net2462[0:1]), .Vd_in_3_col_0(net2466[0:1]), .Vd_in_4_col_0(net2455[0:1]), .Vd_in_5_col_0(net2459[0:1]), .Vd_in_6_col_0(net2463[0:1]), .Vd_in_7_col_0(net2467[0:1]), .Vd_o_0_col_5(net1902[0:1]), .Vd_o_1_col_5(net1903[0:1]), .Vd_o_2_col_5(net1904[0:1]), .Vd_o_3_col_5(net1905[0:1]), .Vd_o_4_col_5(net1906[0:1]), .Vd_o_5_col_5(net1907[0:1]), .Vd_o_6_col_5(net1908[0:1]), .Vd_o_7_col_5(net1909[0:1]));

 	/*Programming Mux */ 


	/* Frame */ 
	tile_analog_frame cab_frame(.pin_layer(METAL3), .N_n_gateEN(net2496), .N_n_programdrain(net2497), .N_n_rundrain(net2498), .N_n_cew0(net2472[0]), .N_n_cew1(net2473[0]), .N_n_cew2(net2474[0]), .N_n_cew3(net2475[0]), .N_n_vtun(net2560[0]), .N_n_vinj_0_(net2503), .N_n_vinj_1_(net2504), .N_n_vinj_2_(net2230[8]), .N_n_gnd_0_(net2505), .N_n_gnd_1_(net2506), .N_n_gnd_2_(net2231[8]), .N_n_avdd(net2507[0]), .N_n_s0(net2476[0]), .N_n_s1(net2477[0]), .N_n_s2(net2478[0]), .N_n_s3(net2479[0]), .N_n_s4(net2480[0]), .N_n_s5(net2481[0]), .N_n_s6(net2482[0]), .N_n_s7(net2483[0]), .N_n_s8(net2484[0]), .N_n_s9(net2485[0]), .N_n_s10(net2486[0]), .N_n_s11(net2487[0]), .N_n_s12(net2488), .N_n_s13(net2489), .N_n_s14(net2490), .N_n_s15(net2491), .N_n_s16(net2492), .N_n_s17(net2493), .N_n_s18(net2494), .N_n_s19(net2495), .N_n_prog(net2528[0]), .N_n_run(net2529), .N_n_vgsel(net2530), .S_s_gateEN(net2496), .S_s_programdrain(net2497), .S_s_rundrain(net2498), .S_s_cew0(net2499[0]), .S_s_cew1(net2500[0]), .S_s_cew2(net2501[0]), .S_s_cew3(net2502[0]), .S_s_vtun(net2560[0]), .S_s_vinj_0_(net2503), .S_s_vinj_1_(net2504), .S_s_vinj_2_(net2230[8]), .S_s_gnd_0_(net2505), .S_s_gnd_1_(net2506), .S_s_gnd_2_(net2231[8]), .S_s_avdd(net2507[0]), .S_s_s0(net2508), .S_s_s1(net2509), .S_s_s2(net2510), .S_s_s3(net2511), .S_s_s4(net2512), .S_s_s5(net2513), .S_s_s6(net2514), .S_s_s7(net2515), .S_s_s8(net2516[0]), .S_s_s9(net2517[0]), .S_s_s10(net2518[0]), .S_s_s11(net2519[0]), .S_s_s12(net2520[0]), .S_s_s13(net2521[0]), .S_s_s14(net2522[0]), .S_s_s15(net2523[0]), .S_s_s16(net2524[0]), .S_s_s17(net2525[0]), .S_s_s18(net2526[0]), .S_s_s19(net2527[0]), .S_s_prog(net2528[0]), .S_s_run(net2529), .S_s_vgsel(net2530), .W_w_cns0(net2499[1]), .W_w_cns1(net2500[1]), .W_w_cns2(net2501[1]), .W_w_cns3(net2502[1]), .W_w_vgrun(net2559[0]), .W_w_vtun(net2560[0]), .W_w_vinj(net2230[8]), .W_w_gnd(net2231[8]), .W_w_avdd(net2563[0]), .W_w_drainbit4(net2564), .W_w_drainbit3(net2565), .W_w_drainbit2(net2566), .W_w_drainbit1(net2567), .W_w_drainbit0(net2568), .W_w_s0(net2535[0]), .W_w_s1(net2536[0]), .W_w_s2(net2537[0]), .W_w_s3(net2538[0]), .W_w_s4(net2539[0]), .W_w_s5(net2540[0]), .W_w_s6(net2541[0]), .W_w_s7(net2542[0]), .W_w_s8(net2543[0]), .W_w_s9(net2544[0]), .W_w_s10(net2545[0]), .W_w_s11(net2546[0]), .W_w_s12(net2547[0]), .W_w_s13(net2548[0]), .W_w_s14(net2549[0]), .W_w_s15(net2550[0]), .W_w_s16(net2551[0]), .W_w_s17(net2552[0]), .W_w_s18(net2553[0]), .W_w_s19(net2554[0]), .W_w_drainbit10(net2589), .W_w_drainbit9(net2590), .W_w_drainbit8(net2591), .W_w_drainbit7(net2592), .W_w_drainbit6(net2593), .W_w_drainbit5(net2594), .W_w_drainEN(net2595), .E_e_cns0(net2555[0]), .E_e_cns1(net2556[0]), .E_e_cns2(net2557[0]), .E_e_cns3(net2558[0]), .E_e_vgrun(net2559[0]), .E_e_vtun(net2560[0]), .E_e_vinj(net2230[8]), .E_e_gnd(net2231[8]), .E_e_avdd(net2563[0]), .E_e_drainbit4(net2564), .E_e_drainbit3(net2565), .E_e_drainbit2(net2566), .E_e_drainbit1(net2567), .E_e_drainbit0(net2568), .E_e_s0(net2569[0]), .E_e_s1(net2570[0]), .E_e_s2(net2571[0]), .E_e_s3(net2572[0]), .E_e_s4(net2569[1]), .E_e_s5(net2570[1]), .E_e_s6(net2571[1]), .E_e_s7(net2572[1]), .E_e_s8(net2569[2]), .E_e_s9(net2570[2]), .E_e_s10(net2571[2]), .E_e_s11(net2572[2]), .E_e_s12(net2569[3]), .E_e_s13(net2570[3]), .E_e_s14(net2571[3]), .E_e_s15(net2572[3]), .E_e_s16(net2569[4]), .E_e_s17(net2570[4]), .E_e_s18(net2571[4]), .E_e_s19(net2572[4]), .E_e_drainbit10(net2589), .E_e_drainbit9(net2590), .E_e_drainbit8(net2591), .E_e_drainbit7(net2592), .E_e_drainbit6(net2593), .E_e_drainbit5(net2594), .E_e_drainEN(net2595));
 endmodule