module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(7), .GND_b_1_row_4(net2221[0:7]), .Vs_b_0_row_4(net124[0:7]), .Vs_b_1_row_4(net125[0:7]), .VINJ_b_1_row_4(net2228[0:7]), .Vsel_b_0_row_4(net2186[0:7]), .Vsel_b_1_row_4(net2187[0:7]), .Vg_b_0_row_4(net2200[0:7]), .Vg_b_1_row_4(net2201[0:7]), .VTUN_brow_4(net2214[0:7]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(17), .matrix_row(5), .matrix_col(9), .GND_b_1_row_4(net2264[0:9]), .Vs_b_0_row_4(net325[0:9]), .Vs_b_1_row_4(net326[0:9]), .VINJ_b_1_row_4(net2263[0:9]), .Vsel_b_0_row_4(net2265[0:9]), .Vsel_b_1_row_4(net2267[0:9]), .Vg_b_0_row_4(net344[0:9]), .Vg_b_1_row_4(net345[0:9]), .VTUN_brow_4(net2262[0:9]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(26), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2241[0:1]), .Vsel_b_0_row_4(net2244[0:1]), .Vsel_b_1_row_4(net2245[0:1]), .Vg_b_0_row_4(net2246[0:1]), .Vg_b_1_row_4(net2247[0:1]), .VTUN_brow_4(net2242[0:1]), .GND_b_1_row_4(net2243[0:1]));
	S_BLOCK_BUFFER I__4 (.island_num(0), .row(0), .col(8), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__5 (.island_num(0), .row(0), .col(9), .matrix_row(4), .matrix_col(1));
	S_BLOCK_CONN_PINS I__6 (.island_num(0), .row(4), .col(9), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__7 (.island_num(0), .row(0), .col(10), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__8 (.island_num(0), .row(3), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__9 (.island_num(0), .row(4), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__10 (.island_num(0), .row(0), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_CONN_PINS I__11 (.island_num(0), .row(2), .col(11), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__12 (.island_num(0), .row(3), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__13 (.island_num(0), .row(0), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_CONN_PINS I__14 (.island_num(0), .row(1), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__15 (.island_num(0), .row(2), .col(12), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__16 (.island_num(0), .row(0), .col(13), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__17 (.island_num(0), .row(1), .col(13), .matrix_row(4), .matrix_col(1));
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2248[0:1]), .Vsel_b_0_row_4(net2251[0:1]), .Vsel_b_1_row_4(net2252[0:1]), .Vg_b_0_row_4(net2253[0:1]), .Vg_b_1_row_4(net2254[0:1]), .VTUN_brow_4(net2249[0:1]), .GND_b_1_row_4(net2250[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2255[0:1]), .Vsel_b_0_row_4(net2258[0:1]), .Vsel_b_1_row_4(net2259[0:1]), .Vg_b_0_row_4(net2260[0:1]), .Vg_b_1_row_4(net2261[0:1]), .VTUN_brow_4(net2256[0:1]), .GND_b_1_row_4(net2257[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(6), .decode_n0_RUN_OUT_0_(net2335), .decode_n0_RUN_OUT_1_(net2336), .decode_n0_RUN_OUT_2_(net2341), .decode_n0_RUN_OUT_3_(net2342), .decode_n1_RUN_OUT_0_(net2347), .decode_n1_RUN_OUT_1_(net2348), .decode_n1_RUN_OUT_2_(net2353), .decode_n1_RUN_OUT_3_(net2354), .decode_n2_RUN_OUT_0_(net2359), .decode_n2_RUN_OUT_1_(net2360), .decode_n2_RUN_OUT_2_(net2365), .decode_n2_RUN_OUT_3_(net2366), .decode_n3_RUN_OUT_0_(net2371), .decode_n3_RUN_OUT_1_(net2372), .decode_n3_RUN_OUT_2_(net2377), .decode_n3_RUN_OUT_3_(net2378), .decode_n4_RUN_OUT_2_(net2383), .decode_n4_RUN_OUT_3_(net2384), .decode_n5_RUN_OUT_0_(net2389), .decode_n5_RUN_OUT_1_(net2390), .decode_n5_RUN_OUT_2_(net2395), .decode_n5_RUN_OUT_3_(net2396), .decode_n6_RUN_OUT_0_(net2401), .decode_n6_RUN_OUT_1_(net2402), .decode_n6_RUN_OUT_2_(net2407), .decode_n6_RUN_OUT_3_(net2408), .decode_n7_RUN_OUT_0_(net2413), .decode_n7_RUN_OUT_1_(net2414), .decode_n7_RUN_OUT_2_(net2419), .decode_n7_RUN_OUT_3_(net2420), .decode_n8_RUN_OUT_0_(net2425), .decode_n8_RUN_OUT_1_(net2426), .decode_n8_RUN_OUT_2_(net2431), .decode_n8_RUN_OUT_3_(net2432), .decode_n9_RUN_OUT_0_(net2437), .decode_n9_RUN_OUT_1_(net2438), .decode_n9_RUN_OUT_2_(net2443), .decode_n9_RUN_OUT_3_(net2444), .decode_n0_OUT_0_(net2333), .decode_n0_OUT_1_(net2334), .decode_n0_OUT_2_(net2339), .decode_n0_OUT_3_(net2340), .decode_n1_OUT_0_(net2345), .decode_n1_OUT_1_(net2346), .decode_n1_OUT_2_(net2351), .decode_n1_OUT_3_(net2352), .decode_n2_OUT_0_(net2357), .decode_n2_OUT_1_(net2358), .decode_n2_OUT_2_(net2363), .decode_n2_OUT_3_(net2364), .decode_n3_OUT_0_(net2369), .decode_n3_OUT_1_(net2370), .decode_n3_OUT_2_(net2375), .decode_n3_OUT_3_(net2376), .decode_n4_OUT_2_(net2381), .decode_n4_OUT_3_(net2382), .decode_n5_OUT_0_(net2387), .decode_n5_OUT_1_(net2388), .decode_n5_OUT_2_(net2393), .decode_n5_OUT_3_(net2394), .decode_n6_OUT_0_(net2399), .decode_n6_OUT_1_(net2400), .decode_n6_OUT_2_(net2405), .decode_n6_OUT_3_(net2406), .decode_n7_OUT_0_(net2411), .decode_n7_OUT_1_(net2412), .decode_n7_OUT_2_(net2417), .decode_n7_OUT_3_(net2418), .decode_n8_OUT_0_(net2423), .decode_n8_OUT_1_(net2424), .decode_n8_OUT_2_(net2429), .decode_n8_OUT_3_(net2430), .decode_n9_OUT_0_(net2435), .decode_n9_OUT_1_(net2436), .decode_n9_OUT_2_(net2441), .decode_n9_OUT_3_(net2442), .decode_n0_VINJ_b_0_(net2331), .decode_n0_VINJ_b_1_(net2337), .decode_n1_VINJ_b_0_(net2343), .decode_n1_VINJ_b_1_(net2349), .decode_n2_VINJ_b_0_(net2355), .decode_n2_VINJ_b_1_(net2361), .decode_n3_VINJ_b_0_(net2367), .decode_n3_VINJ_b_1_(net2373), .decode_n4_VINJ_b_1_(net2379), .decode_n5_VINJ_b_0_(net2385), .decode_n5_VINJ_b_1_(net2391), .decode_n6_VINJ_b_0_(net2397), .decode_n6_VINJ_b_1_(net2403), .decode_n7_VINJ_b_0_(net2409), .decode_n7_VINJ_b_1_(net2415), .decode_n8_VINJ_b_0_(net2421), .decode_n8_VINJ_b_1_(net2427), .decode_n9_VINJ_b_0_(net2433), .decode_n9_VINJ_b_1_(net2439), .decode_n0_GND_b_0_(net2332), .decode_n0_GND_b_1_(net2338), .decode_n1_GND_b_0_(net2344), .decode_n1_GND_b_1_(net2350), .decode_n2_GND_b_0_(net2356), .decode_n2_GND_b_1_(net2362), .decode_n3_GND_b_0_(net2368), .decode_n3_GND_b_1_(net2374), .decode_n4_GND_b_1_(net2380), .decode_n5_GND_b_0_(net2386), .decode_n5_GND_b_1_(net2392), .decode_n6_GND_b_0_(net2398), .decode_n6_GND_b_1_(net2404), .decode_n7_GND_b_0_(net2410), .decode_n7_GND_b_1_(net2416), .decode_n8_GND_b_0_(net2422), .decode_n8_GND_b_1_(net2428), .decode_n9_GND_b_0_(net2434), .decode_n9_GND_b_1_(net2440));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(26), .switch_n0_VPWR_0_(net2335), .switch_n0_VPWR_1_(net2336), .switch_n1_VPWR_0_(net2341), .switch_n1_VPWR_1_(net2342), .switch_n2_VPWR_0_(net2347), .switch_n2_VPWR_1_(net2348), .switch_n3_VPWR_0_(net2353), .switch_n3_VPWR_1_(net2354), .switch_n4_VPWR_0_(net2359), .switch_n4_VPWR_1_(net2360), .switch_n5_VPWR_0_(net2365), .switch_n5_VPWR_1_(net2366), .switch_n6_VPWR_0_(net2371), .switch_n6_VPWR_1_(net2372), .switch_n7_VPWR_0_(net2377), .switch_n7_VPWR_1_(net2378), .switch_n14_VPWR_0_(net2383), .switch_n14_VPWR_1_(net2384), .switch_n16_VPWR_0_(net2389), .switch_n16_VPWR_1_(net2390), .switch_n17_VPWR_0_(net2395), .switch_n17_VPWR_1_(net2396), .switch_n18_VPWR_0_(net2401), .switch_n18_VPWR_1_(net2402), .switch_n19_VPWR_0_(net2407), .switch_n19_VPWR_1_(net2408), .switch_n20_VPWR_0_(net2413), .switch_n20_VPWR_1_(net2414), .switch_n21_VPWR_0_(net2419), .switch_n21_VPWR_1_(net2420), .switch_n22_VPWR_0_(net2425), .switch_n22_VPWR_1_(net2426), .switch_n23_VPWR_0_(net2431), .switch_n23_VPWR_1_(net2432), .switch_n24_VPWR_0_(net2437), .switch_n24_VPWR_1_(net2438), .switch_n25_VPWR_0_(net2443), .switch_n25_VPWR_1_(net2444), .switch_n0_GND_T(net2332), .switch_n1_GND_T(net2338), .switch_n2_GND_T(net2344), .switch_n3_GND_T(net2350), .switch_n4_GND_T(net2356), .switch_n5_GND_T(net2362), .switch_n6_GND_T(net2368), .switch_n7_GND_T(net2374), .switch_n14_GND_T(net2380), .switch_n16_GND_T(net2386), .switch_n17_GND_T(net2392), .switch_n18_GND_T(net2398), .switch_n19_GND_T(net2404), .switch_n20_GND_T(net2410), .switch_n21_GND_T(net2416), .switch_n22_GND_T(net2422), .switch_n23_GND_T(net2428), .switch_n24_GND_T(net2434), .switch_n25_GND_T(net2440), .switch_n0_decode_0_(net2333), .switch_n0_decode_1_(net2334), .switch_n1_decode_0_(net2339), .switch_n1_decode_1_(net2340), .switch_n2_decode_0_(net2345), .switch_n2_decode_1_(net2346), .switch_n3_decode_0_(net2351), .switch_n3_decode_1_(net2352), .switch_n4_decode_0_(net2357), .switch_n4_decode_1_(net2358), .switch_n5_decode_0_(net2363), .switch_n5_decode_1_(net2364), .switch_n6_decode_0_(net2369), .switch_n6_decode_1_(net2370), .switch_n7_decode_0_(net2375), .switch_n7_decode_1_(net2376), .switch_n14_decode_0_(net2381), .switch_n14_decode_1_(net2382), .switch_n16_decode_0_(net2387), .switch_n16_decode_1_(net2388), .switch_n17_decode_0_(net2393), .switch_n17_decode_1_(net2394), .switch_n18_decode_0_(net2399), .switch_n18_decode_1_(net2400), .switch_n19_decode_0_(net2405), .switch_n19_decode_1_(net2406), .switch_n20_decode_0_(net2411), .switch_n20_decode_1_(net2412), .switch_n21_decode_0_(net2417), .switch_n21_decode_1_(net2418), .switch_n22_decode_0_(net2423), .switch_n22_decode_1_(net2424), .switch_n23_decode_0_(net2429), .switch_n23_decode_1_(net2430), .switch_n24_decode_0_(net2435), .switch_n24_decode_1_(net2436), .switch_n25_decode_0_(net2441), .switch_n25_decode_1_(net2442), .switch_n0_VINJ_T(net2331), .switch_n1_VINJ_T(net2337), .switch_n2_VINJ_T(net2343), .switch_n3_VINJ_T(net2349), .switch_n4_VINJ_T(net2355), .switch_n5_VINJ_T(net2361), .switch_n6_VINJ_T(net2367), .switch_n7_VINJ_T(net2373), .switch_n14_VINJ_T(net2379), .switch_n16_VINJ_T(net2385), .switch_n17_VINJ_T(net2391), .switch_n18_VINJ_T(net2397), .switch_n19_VINJ_T(net2403), .switch_n20_VINJ_T(net2409), .switch_n21_VINJ_T(net2415), .switch_n22_VINJ_T(net2421), .switch_n23_VINJ_T(net2427), .switch_n24_VINJ_T(net2433), .switch_n25_VINJ_T(net2439));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch));
	none switch_ind(.island_num(0), .direction(horizontal), .col(8));
	none switch_ind(.island_num(0), .direction(horizontal), .col(9));
	none switch_ind(.island_num(0), .direction(horizontal), .col(10));
	none switch_ind(.island_num(0), .direction(horizontal), .col(11));
	none switch_ind(.island_num(0), .direction(horizontal), .col(12));
	none switch_ind(.island_num(0), .direction(horizontal), .col(13));
	none switch_ind(.island_num(0), .direction(horizontal), .col(15));


	/* Island 1 */
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__0 (.island_num(1), .row(0), .col(0), .matrix_row(1), .matrix_col(8));
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(7), .matrix_col(8), .GND_b_0_row_6(net1223[0:8]), .GND_b_1_row_6(net1224[0:8]), .Vs_b_0_row_6(net1233[0:8]), .Vs_b_1_row_6(net1234[0:8]), .VINJ_b_0_row_6(net1237[0:8]), .VINJ_b_1_row_6(net1238[0:8]), .Vsel_b_0_row_6(net1241[0:8]), .Vsel_b_1_row_6(net1242[0:8]), .Vg_b_0_row_6(net1245[0:8]), .Vg_b_1_row_6(net1246[0:8]), .VTUN_brow_6(net1249[0:8]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(8), .matrix_row(6), .matrix_col(10));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(7), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2086), .P_1_row_0(net2087), .A_0_row_0(net2088), .A_1_row_0(net2089), .A_2_row_0(net2090), .A_3_row_0(net2091));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2099), .P_1_row_0(net2100), .A_0_row_0(net2101), .A_1_row_0(net2102), .A_2_row_0(net2103), .A_3_row_0(net2104));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2117), .P_1_row_0(net2118), .A_0_row_0(net2119), .A_1_row_0(net2120), .A_2_row_0(net2121), .A_3_row_0(net2122));
	TSMC350nm_4TGate_ST_BMatrix_NoSwitch I__8 (.island_num(1), .row(3), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2135), .P_1_row_0(net2136), .P_2_row_0(net2137), .P_3_row_0(net2138), .A_0_row_0(net2139), .A_1_row_0(net2140), .A_2_row_0(net2141), .A_3_row_0(net2142));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2154), .P_1_row_0(net2155), .P_2_row_0(net2156), .P_3_row_0(net2157), .A_0_row_0(net2158), .A_1_row_0(net2159));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net2169), .A_1_row_0(net2170), .A_2_row_0(net2171), .A_3_row_0(net2172));
	TSMC350nm_4TGate_ST_BMatrix I__11 (.island_num(1), .row(6), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net2176), .A_1_row_0(net2177), .A_2_row_0(net2178), .A_3_row_0(net2179));
	TSMC350nm_4TGate_ST_BMatrix I__12 (.island_num(1), .row(7), .col(18), .matrix_row(1), .matrix_col(1));
	TSMC350nm_OutMtrx_IndrctSwcs I__13 (.island_num(1), .row(9), .col(8), .matrix_row(1), .matrix_col(10), .AVDD_rcol_9(net2524[0:1]), .prog_rcol_9(net2525[0:1]));
	TSMC350nm_4x2_Indirect I__14 (.island_num(1), .row(10), .col(8), .matrix_row(2), .matrix_col(10), .Vd_Rl_0_col_0(net1917[0:2]), .Vd_Rl_1_col_0(net1918[0:2]), .Vd_Rl_2_col_0(net1919[0:2]), .Vd_Rl_3_col_0(net1920[0:2]), .Vd_Pl_0_col_0(net1921[0:2]), .Vd_Pl_1_col_0(net1922[0:2]), .Vd_Pl_2_col_0(net1923[0:2]), .Vd_Pl_3_col_0(net1924[0:2]));
	TSMC350nm_4TGate_ST_BMatrix I__15 (.island_num(1), .row(10), .col(18), .matrix_row(2), .matrix_col(1));
	TSMC350nm_TA2Cell_Weak cab_device_16 (.island_num(1), .row(2), .col(19), .VD_P_0_(net2086), .VD_P_1_(net2087), .VIN1_PLUS(net2088), .VIN1_MINUS(net2089), .VIN2_PLUS(net2090), .VIN2_MINUS(net2091), .OUTPUT_0_(net2092[0]), .OUTPUT_1_(net2093[0]), .Vsel_0_(net2163), .Vsel_1_(net2164), .RUN(net2094), .Vg_0_(net2165), .Vg_1_(net2166), .PROG(net2095), .VTUN(net2096), .VINJ(net2097), .GND(net2098), .VPWR(net2524[0]), .Vsel_b_0_(net2107), .Vsel_b_1_(net2108), .RUN_b(net2109), .Vg_b_0_(net2110), .Vg_b_1_(net2111), .PROG_b(net2112), .VTUN_b(net2113), .VINJ_b(net2114), .GND_b(net2115), .VPWR_b(net2116));
	TSMC350nm_TA2Cell_Weak cab_device_17 (.island_num(1), .row(3), .col(19), .VD_P_0_(net2099), .VD_P_1_(net2100), .VIN1_PLUS(net2101), .VIN1_MINUS(net2102), .VIN2_PLUS(net2103), .VIN2_MINUS(net2104), .OUTPUT_0_(net2105[0]), .OUTPUT_1_(net2106[0]), .Vsel_0_(net2107), .Vsel_1_(net2108), .RUN(net2109), .Vg_0_(net2110), .Vg_1_(net2111), .PROG(net2112), .VTUN(net2113), .VINJ(net2114), .GND(net2115), .VPWR(net2116), .Vsel_b_0_(net2125), .Vsel_b_1_(net2126), .RUN_b(net2127), .Vg_b_0_(net2128), .Vg_b_1_(net2129), .PROG_b(net2130), .VTUN_b(net2131), .VINJ_b(net2132), .GND_b(net2133), .VPWR_b(net2134));
	TSMC350nm_TA2Cell_Strong cab_device_18 (.island_num(1), .row(4), .col(19), .VD_P_0_(net2117), .VD_P_1_(net2118), .VIN1_PLUS(net2119), .VIN1_MINUS(net2120), .VIN2_PLUS(net2121), .VIN2_MINUS(net2122), .OUTPUT_0_(net2123[0]), .OUTPUT_1_(net2124[0]), .Vsel_0_(net2125), .Vsel_1_(net2126), .RUN(net2127), .Vg_0_(net2128), .Vg_1_(net2129), .PROG(net2130), .VTUN(net2131), .VINJ(net2132), .GND(net2133), .VPWR(net2134), .Vg_b_0_(net2150), .PROG_b(net2153), .VTUN_b(net2151), .VINJ_b(net2149), .GND_b(net2152));
	TSMC350nm_4WTA_IndirectProg cab_device_19 (.island_num(1), .row(5), .col(19), .VD_P_0_(net2135), .VD_P_1_(net2136), .VD_P_2_(net2137), .VD_P_3_(net2138), .Iin_0_(net2139), .Iin_1_(net2140), .Iin_2_(net2141), .Iin_3_(net2142), .Vout_0_(net2143[0]), .Vout_1_(net2144[0]), .Vout_2_(net2145[0]), .Vout_3_(net2146[0]), .Vmid(net2147[0]), .Vbias(net2148[0]), .Vsel(net2163), .Vs(net2524[0]), .VINJ(net2149), .Vg(net2150), .VTUN(net2151), .GND(net2152), .PROG(net2153), .VINJ_b(net2162), .VTUN_b(net2168), .GND_b(net2167));
	TSMC350nm_Cap_Bank cab_device_20 (.island_num(1), .row(6), .col(19), .VD_P_0_(net2154), .VD_P_1_(net2155), .VD_P_2_(net2156), .VD_P_3_(net2157), .VIN_0_(net2158), .VIN_1_(net2159), .OUT_0_(net2160[0]), .OUT_1_(net2161[0]), .VINJ(net2162), .Vsel_0_(net2163), .Vsel_1_(net2164), .Vg_0_(net2165), .Vg_1_(net2166), .GND(net2167), .VTUN(net2168), .GND_b(net2175));
	TSMC350nm_NandPfets cab_device_21 (.island_num(1), .row(7), .col(19), .GATE_N(net2169), .SOURCE_N(net2170), .GATE_P(net2171), .SOURCE_P(net2172), .DRAIN_N(net2173[0]), .DRAIN_P(net2174[0]), .VPWR(net2524[0]), .GND(net2175), .VPWR_b(net2183), .GND_b(net2184));
	TSMC350nm_TGate_2nMirror cab_device_22 (.island_num(1), .row(8), .col(19), .IN_CM_0_(net2176), .IN_CM_1_(net2177), .SelN(net2178), .IN_TG(net2179), .OUT_CM_0_(net2180[0]), .OUT_CM_1_(net2181[0]), .OUT_TG(net2182[0]), .VPWR(net2183), .GND(net2184));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(1), .direction(vertical), .num(12), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(12), .type(prog_switch), .switch_n8_PR_0_(net2509[0]), .switch_n8_PR_1_(net2513[0]), .switch_n8_PR_2_(net2517[0]), .switch_n8_PR_3_(net2521[0]), .switch_n8_In_0_(net2508[0]), .switch_n8_In_1_(net2512[0]), .switch_n8_In_2_(net2516[0]), .switch_n8_In_3_(net2520[0]));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(20), .switch_n0_Input_0_(net2185), .switch_n0_Input_1_(net2221[0]), .switch_n1_Input_0_(net124[1]), .switch_n1_Input_1_(net125[1]), .switch_n2_Input_0_(net124[2]), .switch_n2_Input_1_(net125[2]), .switch_n3_Input_0_(net124[3]), .switch_n3_Input_1_(net125[3]), .switch_n4_Input_0_(net325[0]), .switch_n4_Input_1_(net326[0]), .switch_n5_Input_0_(net325[1]), .switch_n5_Input_1_(net326[1]), .switch_n6_Input_0_(net325[2]), .switch_n6_Input_1_(net326[2]), .switch_n7_Input_0_(net325[3]), .switch_n7_Input_1_(net326[3]), .switch_n8_Input_0_(net2507[0]), .switch_n8_Input_1_(net2092[0]), .switch_n9_Input_0_(net2093[0]), .switch_n9_Input_1_(net2105[0]), .switch_n10_Input_0_(net2106[0]), .switch_n10_Input_1_(net2123[0]), .switch_n11_Input_0_(net2124[0]), .switch_n11_Input_1_(net2143[0]), .switch_n12_Input_0_(net2144[0]), .switch_n12_Input_1_(net2145[0]), .switch_n13_Input_0_(net2146[0]), .switch_n13_Input_1_(net2147[0]), .switch_n14_Input_0_(net2148[0]), .switch_n14_Input_1_(net2160[0]), .switch_n15_Input_0_(net2161[0]), .switch_n15_Input_1_(net2173[0]), .switch_n16_Input_0_(net2174[0]), .switch_n16_Input_1_(net2180[0]), .switch_n17_Input_0_(net2181[0]), .switch_n17_Input_1_(net2182[0]), .switch_n0_GND(net2221[0]), .switch_n1_GND(net2221[1]), .switch_n2_GND(net2221[2]), .switch_n3_GND(net2221[3]), .switch_n4_GND(net2221[4]), .switch_n5_GND(net2221[5]), .switch_n6_GND(net2221[6]), .switch_n7_GND(net2243[0]), .switch_n8_GND(net2250[0]), .switch_n9_GND(net2257[0]), .switch_n10_GND(net2264[0]), .switch_n11_GND(net2264[1]), .switch_n12_GND(net2264[2]), .switch_n13_GND(net2264[3]), .switch_n14_GND(net2264[4]), .switch_n15_GND(net2264[5]), .switch_n16_GND(net2264[6]), .switch_n17_GND(net2264[7]), .switch_n0_Vsel_0_(net2186[0]), .switch_n0_Vsel_1_(net2187[0]), .switch_n1_Vsel_0_(net2186[1]), .switch_n1_Vsel_1_(net2187[1]), .switch_n2_Vsel_0_(net2186[2]), .switch_n2_Vsel_1_(net2187[2]), .switch_n3_Vsel_0_(net2186[3]), .switch_n3_Vsel_1_(net2187[3]), .switch_n4_Vsel_0_(net2186[4]), .switch_n4_Vsel_1_(net2187[4]), .switch_n5_Vsel_0_(net2186[5]), .switch_n5_Vsel_1_(net2187[5]), .switch_n6_Vsel_0_(net2186[6]), .switch_n6_Vsel_1_(net2187[6]), .switch_n7_Vsel_0_(net2245[0]), .switch_n7_Vsel_1_(net2244[0]), .switch_n8_Vsel_0_(net2252[0]), .switch_n8_Vsel_1_(net2251[0]), .switch_n9_Vsel_0_(net2259[0]), .switch_n9_Vsel_1_(net2258[0]), .switch_n10_Vsel_0_(net2265[0]), .switch_n10_Vsel_1_(net2267[0]), .switch_n11_Vsel_0_(net2265[1]), .switch_n11_Vsel_1_(net2267[1]), .switch_n12_Vsel_0_(net2265[2]), .switch_n12_Vsel_1_(net2267[2]), .switch_n13_Vsel_0_(net2265[3]), .switch_n13_Vsel_1_(net2267[3]), .switch_n14_Vsel_0_(net2265[4]), .switch_n14_Vsel_1_(net2267[4]), .switch_n15_Vsel_0_(net2265[5]), .switch_n15_Vsel_1_(net2267[5]), .switch_n16_Vsel_0_(net2265[6]), .switch_n16_Vsel_1_(net2267[6]), .switch_n17_Vsel_0_(net2265[7]), .switch_n17_Vsel_1_(net2267[7]), .switch_n0_Vg_global_0_(net2200[0]), .switch_n0_Vg_global_1_(net2201[0]), .switch_n1_Vg_global_0_(net2200[1]), .switch_n1_Vg_global_1_(net2201[1]), .switch_n2_Vg_global_0_(net2200[2]), .switch_n2_Vg_global_1_(net2201[2]), .switch_n3_Vg_global_0_(net2200[3]), .switch_n3_Vg_global_1_(net2201[3]), .switch_n4_Vg_global_0_(net2200[4]), .switch_n4_Vg_global_1_(net2201[4]), .switch_n5_Vg_global_0_(net2200[5]), .switch_n5_Vg_global_1_(net2201[5]), .switch_n6_Vg_global_0_(net2200[6]), .switch_n6_Vg_global_1_(net2201[6]), .switch_n7_Vg_global_0_(net2247[0]), .switch_n7_Vg_global_1_(net2246[0]), .switch_n8_Vg_global_0_(net2254[0]), .switch_n8_Vg_global_1_(net2253[0]), .switch_n9_Vg_global_0_(net2261[0]), .switch_n9_Vg_global_1_(net2260[0]), .switch_n10_Vg_global_0_(net344[0]), .switch_n10_Vg_global_1_(net345[0]), .switch_n11_Vg_global_0_(net344[1]), .switch_n11_Vg_global_1_(net345[1]), .switch_n12_Vg_global_0_(net344[2]), .switch_n12_Vg_global_1_(net345[2]), .switch_n13_Vg_global_0_(net344[3]), .switch_n13_Vg_global_1_(net345[3]), .switch_n14_Vg_global_0_(net344[4]), .switch_n14_Vg_global_1_(net345[4]), .switch_n15_Vg_global_0_(net344[5]), .switch_n15_Vg_global_1_(net345[5]), .switch_n16_Vg_global_0_(net344[6]), .switch_n16_Vg_global_1_(net345[6]), .switch_n17_Vg_global_0_(net344[7]), .switch_n17_Vg_global_1_(net345[7]), .switch_n0_VTUN(net2214[0]), .switch_n1_VTUN(net2214[1]), .switch_n2_VTUN(net2214[2]), .switch_n3_VTUN(net2214[3]), .switch_n4_VTUN(net2214[4]), .switch_n5_VTUN(net2214[5]), .switch_n6_VTUN(net2214[6]), .switch_n7_VTUN(net2242[0]), .switch_n8_VTUN(net2249[0]), .switch_n9_VTUN(net2256[0]), .switch_n10_VTUN(net2262[0]), .switch_n11_VTUN(net2262[1]), .switch_n12_VTUN(net2262[2]), .switch_n13_VTUN(net2262[3]), .switch_n14_VTUN(net2262[4]), .switch_n15_VTUN(net2262[5]), .switch_n16_VTUN(net2262[6]), .switch_n17_VTUN(net2262[7]), .switch_n0_VINJ(net2228[0]), .switch_n1_VINJ(net2228[1]), .switch_n2_VINJ(net2228[2]), .switch_n3_VINJ(net2228[3]), .switch_n4_VINJ(net2228[4]), .switch_n5_VINJ(net2228[5]), .switch_n6_VINJ(net2228[6]), .switch_n7_VINJ(net2241[0]), .switch_n8_VINJ(net2248[0]), .switch_n9_VINJ(net2255[0]), .switch_n10_VINJ(net2263[0]), .switch_n11_VINJ(net2263[1]), .switch_n12_VINJ(net2263[2]), .switch_n13_VINJ(net2263[3]), .switch_n14_VINJ(net2263[4]), .switch_n15_VINJ(net2263[5]), .switch_n16_VINJ(net2263[6]), .switch_n17_VINJ(net2263[7]), .switch_n0_AVDD_r(net2524[0]));
	none switch_ind(.island_num(1), .direction(horizontal), .col(18));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(19), .VPWR_0_(net2185), .VPWR_1_(net2185), .GND_T(net2264[8]), .VTUN_T(net2262[8]), .decode_0_(net2265[8]), .decode_1_(net2267[8]), .VINJ_T(net2263[8]), .GND(net2098), .CTRL_B_0_(net2163), .CTRL_B_1_(net2164), .run_r(net2094), .prog_r(net2095), .Vg_0_(net2165), .Vg_1_(net2166), .VTUN(net2096), .VINJ(net2097), .VDD_1_(net2524[0]), .PROG(net2525[0]));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net1233[0:6]), .out_1_row_0(net1234[0:6]), .VINJ_0_row_0(net1237[0:6]), .VINJ_1_row_0(net1238[0:6]), .Vsel_0_row_0(net1241[0:6]), .Vsel_1_row_0(net1242[0:6]), .Vg_0_row_0(net1245[0:6]), .Vg_1_row_0(net1246[0:6]), .GNDrow_0(net1223[0:6]), .VTUNrow_0(net1249[0:6]), .Dcol_0(net124[6:7]), .CLKcol_0(net125[6:7]), .Qcol_5(net125[6:7]), .comcol_0(net2507[0:1]), .VDDcol_0(net2524[0:1]), .Vd_Pcol_0(net2521[0:1]), .Vd_in_0_col_0(net2508[0:1]), .Vd_in_1_col_0(net2512[0:1]), .Vd_in_2_col_0(net2516[0:1]), .Vd_in_3_col_0(net2520[0:1]), .Vd_in_4_col_0(net2509[0:1]), .Vd_in_5_col_0(net2513[0:1]), .Vd_in_6_col_0(net2517[0:1]), .Vd_in_7_col_0(net2521[0:1]), .Vd_o_0_col_5(net1917[0:1]), .Vd_o_1_col_5(net1918[0:1]), .Vd_o_2_col_5(net1919[0:1]), .Vd_o_3_col_5(net1920[0:1]), .Vd_o_4_col_5(net1921[0:1]), .Vd_o_5_col_5(net1922[0:1]), .Vd_o_6_col_5(net1923[0:1]), .Vd_o_7_col_5(net1924[0:1]));

 	/*Programming Mux */ 

 endmodule