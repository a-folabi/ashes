module cells_only(port1);

ArbGen I__0 (.island_num(0), .row(1), .col(1), .Vout_0_(net0), .Vout_1_(net1), .Vout_2_(net2), .Vout_3_(net3), .Vout_4_(net4), .Vout_5_(net5), .Vout_6_(net6), .Vout_7_(net7), .Vout_8_(net8), .Vout_9_(net9), .Vout_10_(net10), .Vout_11_(net11), .Vout_12_(net12), .Vout_13_(net13), .Vout_14_(net14), .Vout_15_(net15), .Vout_16_(net16), .Vout_17_(net17), .Vout_18_(net18), .Vout_19_(net19), .Vout_20_(net20), .Vout_21_(net21), .Vout_22_(net22), .Vout_23_(net23), .Vout_24_(net24), .Vout_25_(net25), .Vout_26_(net26), .Vout_27_(net27), .Vout_28_(net28), .Vout_29_(net29), .Vout_30_(net30), .Vout_31_(net31), .Vout_32_(net32), .Vout_33_(net33), .Vout_34_(net34), .Vout_35_(net35), .Vout_36_(net36), .Vout_37_(net37), .Vout_38_(net38), .Vout_39_(net39), .Vout_40_(net40), .Vout_41_(net41), .Vout_42_(net42), .Vout_43_(net43), .Vout_44_(net44), .Vout_45_(net45), .Vout_46_(net46), .Vout_47_(net47), .Vout_48_(net48), .Vout_49_(net49), .Vout_50_(net50), .Vout_51_(net51), .Vout_52_(net52), .Vout_53_(net53), .Vout_54_(net54), .Vout_55_(net55), .Vout_56_(net56), .Vout_57_(net57), .Vout_58_(net58), .Vout_59_(net59), .Vout_60_(net60), .Vout_61_(net61), .Vout_62_(net62), .Vout_63_(net63));

Classifer_64x64 I__1 (.island_num(1), .row(1), .col(1), .VGRUN_0_(net0), .VGRUN_1_(net1), .VGRUN_2_(net2), .VGRUN_3_(net3), .VGRUN_4_(net4), .VGRUN_5_(net5), .VGRUN_6_(net6), .VGRUN_7_(net7), .VGRUN_8_(net8), .VGRUN_9_(net9), .VGRUN_10_(net10), .VGRUN_11_(net11), .VGRUN_12_(net12), .VGRUN_13_(net13), .VGRUN_14_(net14), .VGRUN_15_(net15), .VGRUN_16_(net16), .VGRUN_17_(net17), .VGRUN_18_(net18), .VGRUN_19_(net19), .VGRUN_20_(net20), .VGRUN_21_(net21), .VGRUN_22_(net22), .VGRUN_23_(net23), .VGRUN_24_(net24), .VGRUN_25_(net25), .VGRUN_26_(net26), .VGRUN_27_(net27), .VGRUN_28_(net28), .VGRUN_29_(net29), .VGRUN_30_(net30), .VGRUN_31_(net31), .VGRUN_32_(net32), .VGRUN_33_(net33), .VGRUN_34_(net34), .VGRUN_35_(net35), .VGRUN_36_(net36), .VGRUN_37_(net37), .VGRUN_38_(net38), .VGRUN_39_(net39), .VGRUN_40_(net40), .VGRUN_41_(net41), .VGRUN_42_(net42), .VGRUN_43_(net43), .VGRUN_44_(net44), .VGRUN_45_(net45), .VGRUN_46_(net46), .VGRUN_47_(net47), .VGRUN_48_(net48), .VGRUN_49_(net49), .VGRUN_50_(net50), .VGRUN_51_(net51), .VGRUN_52_(net52), .VGRUN_53_(net53), .VGRUN_54_(net54), .VGRUN_55_(net55), .VGRUN_56_(net56), .VGRUN_57_(net57), .VGRUN_58_(net58), .VGRUN_59_(net59), .VGRUN_60_(net60), .VGRUN_61_(net61), .VGRUN_62_(net62), .VGRUN_63_(net63), .OUT_0_(net64), .OUT_1_(net65), .OUT_2_(net66), .OUT_3_(net67), .OUT_4_(net68), .OUT_5_(net69), .OUT_6_(net70), .OUT_7_(net71), .OUT_8_(net72), .OUT_9_(net73), .OUT_10_(net74), .OUT_11_(net75), .OUT_12_(net76), .OUT_13_(net77), .OUT_14_(net78), .OUT_15_(net79), .OUT_16_(net80), .OUT_17_(net81), .OUT_18_(net82), .OUT_19_(net83), .OUT_20_(net84), .OUT_21_(net85), .OUT_22_(net86), .OUT_23_(net87), .OUT_24_(net88), .OUT_25_(net89), .OUT_26_(net90), .OUT_27_(net91), .OUT_28_(net92), .OUT_29_(net93), .OUT_30_(net94), .OUT_31_(net95), .OUT_32_(net96), .OUT_33_(net97), .OUT_34_(net98), .OUT_35_(net99), .OUT_36_(net100), .OUT_37_(net101), .OUT_38_(net102), .OUT_39_(net103), .OUT_40_(net104), .OUT_41_(net105), .OUT_42_(net106), .OUT_43_(net107), .OUT_44_(net108), .OUT_45_(net109), .OUT_46_(net110), .OUT_47_(net111), .OUT_48_(net112), .OUT_49_(net113), .OUT_50_(net114), .OUT_51_(net115), .OUT_52_(net116), .OUT_53_(net117), .OUT_54_(net118), .OUT_55_(net119), .OUT_56_(net120), .OUT_57_(net121), .OUT_58_(net122), .OUT_59_(net123), .OUT_60_(net124), .OUT_61_(net125), .OUT_62_(net126), .OUT_63_(net127));

SpeedTest_DigitalReadout_64x32 I__2 (.island_num(2), .row(1), .col(1), .Din_0_(net64), .Din_1_(net65), .Din_2_(net66), .Din_3_(net67), .Din_4_(net68), .Din_5_(net69), .Din_6_(net70), .Din_7_(net71), .Din_8_(net72), .Din_9_(net73), .Din_10_(net74), .Din_11_(net75), .Din_12_(net76), .Din_13_(net77), .Din_14_(net78), .Din_15_(net79), .Din_16_(net80), .Din_17_(net81), .Din_18_(net82), .Din_19_(net83), .Din_20_(net84), .Din_21_(net85), .Din_22_(net86), .Din_23_(net87), .Din_24_(net88), .Din_25_(net89), .Din_26_(net90), .Din_27_(net91), .Din_28_(net92), .Din_29_(net93), .Din_30_(net94), .Din_31_(net95), .Din_32_(net96), .Din_33_(net97), .Din_34_(net98), .Din_35_(net99), .Din_36_(net100), .Din_37_(net101), .Din_38_(net102), .Din_39_(net103), .Din_40_(net104), .Din_41_(net105), .Din_42_(net106), .Din_43_(net107), .Din_44_(net108), .Din_45_(net109), .Din_46_(net110), .Din_47_(net111), .Din_48_(net112), .Din_49_(net113), .Din_50_(net114), .Din_51_(net115), .Din_52_(net116), .Din_53_(net117), .Din_54_(net118), .Din_55_(net119), .Din_56_(net120), .Din_57_(net121), .Din_58_(net122), .Din_59_(net123), .Din_60_(net124), .Din_61_(net125), .Din_62_(net126), .Din_63_(net127));

endmodule