module TOP(port1);


	/* Island 0 */
	TSMC350nm_C4 I__0 (.island_num(0), .row(0), .col(0), .matrix_row(12), .matrix_col(1), .OUTPUTcol_0(net232[0:12]));

 	/*Programming Mux */ 


	/* Island 1 */
	TSMC350nm_Ampdet_NoFG I__0 (.island_num(1), .row(0), .col(0), .matrix_row(12), .matrix_col(1), .VINcol_0(net232[0:12]), .OUTPUTcol_0(net244[0:12]));

 	/*Programming Mux */ 


	/* Island 2 */
	TSMC350nm_DelayBlock_3stage_new I__0 (.island_num(2), .row(0), .col(0), .matrix_row(12), .matrix_col(1), .VINcol_0(net244[0:12]), .VOUT_0_col_0(net611[0:12]), .VOUT_1_col_0(net612[0:12]), .VOUT_2_col_0(net613[0:12]));

 	/*Programming Mux */ 


	/* Island 3 */
	TSMC350nm_VMMWTA I__0 (.island_num(3), .row(0), .col(17), .matrix_row(9), .matrix_col(1), .matrix_row(9), .matrix_col(1));
	TSMC350nm_4x2_Indirect I__1 (.island_num(3), .row(0), .col(0), .matrix_row(9), .matrix_col(17));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(3), .direction(horizontal), .bits(6), .decode_n0_VGRUN_0_(net611[0]), .decode_n0_VGRUN_1_(net612[0]), .decode_n0_VGRUN_2_(net613[0]), .decode_n0_VGRUN_3_(net614[0]), .decode_n1_VGRUN_0_(net611[1]), .decode_n1_VGRUN_1_(net612[1]), .decode_n1_VGRUN_2_(net613[1]), .decode_n1_VGRUN_3_(net614[1]), .decode_n2_VGRUN_0_(net611[2]), .decode_n2_VGRUN_1_(net612[2]), .decode_n2_VGRUN_2_(net613[2]), .decode_n2_VGRUN_3_(net614[2]), .decode_n3_VGRUN_0_(net611[3]), .decode_n3_VGRUN_1_(net612[3]), .decode_n3_VGRUN_2_(net613[3]), .decode_n3_VGRUN_3_(net614[3]), .decode_n4_VGRUN_0_(net611[4]), .decode_n4_VGRUN_1_(net612[4]), .decode_n4_VGRUN_2_(net613[4]), .decode_n4_VGRUN_3_(net614[4]), .decode_n5_VGRUN_0_(net611[5]), .decode_n5_VGRUN_1_(net612[5]), .decode_n5_VGRUN_2_(net613[5]), .decode_n5_VGRUN_3_(net614[5]), .decode_n6_VGRUN_0_(net611[6]), .decode_n6_VGRUN_1_(net612[6]), .decode_n6_VGRUN_2_(net613[6]), .decode_n6_VGRUN_3_(net614[6]), .decode_n7_VGRUN_0_(net611[7]), .decode_n7_VGRUN_1_(net612[7]), .decode_n7_VGRUN_2_(net613[7]), .decode_n7_VGRUN_3_(net614[7]), .decode_n8_VGRUN_0_(net611[8]), .decode_n8_VGRUN_1_(net612[8]), .decode_n8_VGRUN_2_(net613[8]), .decode_n8_VGRUN_3_(net614[8]));
	TSMC350nm_IndirectSwitches switch(.island_num(3), .direction(horizontal), .num(18));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(3), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect01d3 switch(.island_num(3), .direction(vertical), .num(9), .type(drain_select));
	TSMC350nm_FourTgate_ThickOx_FG_MEM switch(.island_num(3), .direction(vertical), .num(9), .type(prog_switch));
endmodule