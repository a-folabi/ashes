VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER routingPitch REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.01 ;
LAYER POLY1
  TYPE MASTERSLICE ;
END POLY1

LAYER CONT
  TYPE CUT ;
  SPACING 0.4 ;
END CONT

LAYER METAL1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.5 ;
  SPACING 0.45 ;
  PROPERTY routingPitch 1.25 ;
END METAL1

LAYER VIA12
  TYPE CUT ;
  SPACING 0.45 ;
END VIA12

LAYER METAL2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.4 ;
END METAL2

LAYER VIA23
  TYPE CUT ;
  SPACING 0.45 ;
END VIA23

LAYER METAL3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.25 ;
END METAL3

LAYER VIA34
  TYPE CUT ;
  SPACING 0.45 ;
END VIA34

LAYER METAL4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.6 ;
  PROPERTY routingPitch 1.4 ;
END METAL4

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIARULE M4_M3 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL4 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1

VIARULE M1_POLY1 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 1 ;
END M1_POLY1

VIA M1_POLY1s
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER POLY1 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.35 -0.35 0.35 0.35 ;
END M1_POLY1s

VIA M2_M1s
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL2 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M2_M1s

VIA M3_M2s
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL3 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL2 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M3_M2s

VIA M4_M3s
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL3 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M4_M3s

VIARULE openMSP430_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END openMSP430_VIA0

VIARULE openMSP430_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END openMSP430_VIA1

VIARULE analog_mem_ctrlr_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END analog_mem_ctrlr_VIA4

VIARULE analog_mem_ctrlr_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END analog_mem_ctrlr_VIA3

VIARULE analog_mem_ctrlr_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END analog_mem_ctrlr_VIA2

VIARULE analog_mem_ctrlr_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END analog_mem_ctrlr_VIA1

VIARULE analog_mem_ctrlr_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END analog_mem_ctrlr_VIA0

VIARULE dacbank_periph_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_periph_VIA0

VIARULE dacbank_periph_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_periph_VIA2

VIARULE dacbank_periph_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_periph_VIA1

VIARULE dacbank_periph_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_periph_VIA3

VIARULE dacbank_periph_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_periph_VIA4

VIARULE dacbank_periph_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_periph_VIA5

VIARULE dacbank_periph_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_periph_VIA7

VIARULE openMSP430_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END openMSP430_VIA2

VIARULE gp_per160_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per160_VIA4

VIARULE gp_per160_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per160_VIA3

VIARULE gp_per160_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per160_VIA2

VIARULE gp_per160_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END gp_per160_VIA1

VIARULE gp_per160_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END gp_per160_VIA0

VIARULE gp_per168_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per168_VIA4

VIARULE gp_per168_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per168_VIA3

VIARULE gp_per168_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per168_VIA2

VIARULE gp_per168_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END gp_per168_VIA1

VIARULE gp_per168_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END gp_per168_VIA0

VIARULE gp_per170_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per170_VIA4

VIARULE gp_per170_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per170_VIA3

VIARULE gp_per170_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per170_VIA2

VIARULE gp_per170_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END gp_per170_VIA1

VIARULE gp_per170_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END gp_per170_VIA0

VIARULE gp_per_in178_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per_in178_VIA4

VIARULE gp_per_in178_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per_in178_VIA3

VIARULE gp_per_in178_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END gp_per_in178_VIA2

VIARULE gp_per_in178_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END gp_per_in178_VIA1

VIARULE gp_per_in178_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END gp_per_in178_VIA0

VIARULE spi_master_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END spi_master_VIA4

VIARULE spi_master_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END spi_master_VIA3

VIARULE spi_master_VIA2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END spi_master_VIA2

VIARULE spi_master_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END spi_master_VIA1

VIARULE spi_master_VIA0 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END spi_master_VIA0

VIARULE spi_periph_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END spi_periph_VIA4

VIARULE spi_periph_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END spi_periph_VIA3

VIARULE spi_periph_VIA2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END spi_periph_VIA2

VIARULE spi_periph_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END spi_periph_VIA1

VIARULE spi_periph_VIA0 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END spi_periph_VIA0

VIARULE memctrlr_cadsp_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END memctrlr_cadsp_VIA7

VIARULE comm_aer_out_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END comm_aer_out_VIA4

VIARULE comm_aer_out_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END comm_aer_out_VIA3

VIARULE comm_aer_out_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END comm_aer_out_VIA2

VIARULE comm_aer_out_VIA1 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END comm_aer_out_VIA1

VIARULE comm_aer_out_VIA0 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END comm_aer_out_VIA0

VIARULE comm_aer_in_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END comm_aer_in_VIA0

VIARULE comm_aer_in_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END comm_aer_in_VIA1

VIARULE comm_aer_in_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END comm_aer_in_VIA2

VIARULE comm_aer_in_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END comm_aer_in_VIA3

VIARULE comm_aer_in_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END comm_aer_in_VIA4

VIARULE aer_in256_lo_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in256_lo_VIA4

VIARULE aer_in256_lo_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in256_lo_VIA3

VIARULE aer_in256_lo_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in256_lo_VIA2

VIARULE aer_in256_lo_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in256_lo_VIA1

VIARULE aer_in256_lo_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in256_lo_VIA0

VIARULE aer_in256_hi_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in256_hi_VIA4

VIARULE aer_in256_hi_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in256_hi_VIA3

VIARULE aer_in256_hi_VIA2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in256_hi_VIA2

VIARULE aer_in256_hi_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in256_hi_VIA1

VIARULE aer_in256_hi_VIA0 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in256_hi_VIA0

VIARULE aer_out256_VIA9 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out256_VIA9

VIARULE aer_out256_VIA8 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out256_VIA8

VIARULE aer_out256_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.475 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.475 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out256_VIA7

VIARULE aer_out256_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.475 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.475 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out256_VIA6

VIARULE aer_out256_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out256_VIA5

VIARULE aer_out256_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out256_VIA4

VIARULE aer_out256_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out256_VIA3

VIARULE aer_out256_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out256_VIA2

VIARULE aer_out256_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_out256_VIA1

VIARULE aer_out256_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_out256_VIA0

VIARULE periph_neuron2_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_neuron2_VIA4

VIARULE periph_neuron2_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_neuron2_VIA3

VIARULE periph_neuron2_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END periph_neuron2_VIA2

VIARULE periph_neuron2_VIA1 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END periph_neuron2_VIA1

VIARULE periph_neuron2_VIA0 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_neuron2_VIA0

VIARULE aer_out70_VIA9 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out70_VIA9

VIARULE aer_out70_VIA8 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out70_VIA8

VIARULE aer_out70_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.475 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.475 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out70_VIA7

VIARULE aer_out70_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.475 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.475 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out70_VIA6

VIARULE aer_out70_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out70_VIA5

VIARULE aer_out70_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out70_VIA4

VIARULE aer_out70_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_out70_VIA3

VIARULE aer_out70_VIA2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_out70_VIA2

VIARULE aer_out70_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out70_VIA1

VIARULE aer_out70_VIA0 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out70_VIA0

VIARULE aer_in200_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in200_VIA4

VIARULE aer_in200_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in200_VIA3

VIARULE aer_in200_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in200_VIA2

VIARULE aer_in200_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in200_VIA1

VIARULE aer_in200_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in200_VIA0

VIARULE periph_1h_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_1h_VIA7

VIARULE periph_1h_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_1h_VIA6

VIARULE periph_1h_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_1h_VIA5

VIARULE periph_1h_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_1h_VIA4

VIARULE periph_1h_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_1h_VIA3

VIARULE periph_1h_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END periph_1h_VIA2

VIARULE periph_1h_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END periph_1h_VIA1

VIARULE periph_1h_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END periph_1h_VIA0

VIARULE dacbank_x12_periph_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END dacbank_x12_periph_VIA0

VIARULE dacbank_x12_periph_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_x12_periph_VIA1

VIARULE dacbank_x12_periph_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_x12_periph_VIA2

VIARULE dacbank_x12_periph_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END dacbank_x12_periph_VIA3

VIARULE dacbank_x12_periph_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_x12_periph_VIA4

VIARULE rain_periph_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END rain_periph_VIA0

VIARULE rain_periph_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END rain_periph_VIA1

VIARULE rain_periph_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END rain_periph_VIA2

VIARULE rain_periph_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END rain_periph_VIA3

VIARULE rain_periph_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.3 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END rain_periph_VIA4

VIARULE aer_out400_VIA0 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out400_VIA0

VIARULE aer_out400_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out400_VIA1

VIARULE aer_out400_VIA2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_out400_VIA2

VIARULE aer_out400_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_out400_VIA3

VIARULE aer_out400_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out400_VIA4

VIARULE aer_out400_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out400_VIA5

VIARULE aer_out400_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.475 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.475 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out400_VIA6

VIARULE aer_out400_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.475 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.475 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out400_VIA7

VIARULE aer_out400_VIA8 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out400_VIA8

VIARULE aer_out400_VIA9 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out400_VIA9

VIARULE aer_in300_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in300_VIA4

VIARULE aer_in300_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in300_VIA3

VIARULE aer_in300_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.35 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in300_VIA2

VIARULE aer_in300_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in300_VIA1

VIARULE aer_in300_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in300_VIA0

VIARULE aer_in300_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in300_VIA5

VIARULE aer_in300_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.475 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.475 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in300_VIA6

VIARULE aer_in300_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.475 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.475 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in300_VIA7

VIARULE aer_in300_VIA8 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.475 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in300_VIA8

VIARULE aer_in300_VIA9 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in300_VIA9

VIARULE aer_out_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_out_VIA0

VIARULE aer_out_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_out_VIA1

VIARULE aer_out_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out_VIA2

VIARULE aer_out_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out_VIA3

VIARULE aer_out_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out_VIA4

VIARULE aer_out_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out_VIA5

VIARULE aer_out_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out_VIA6

VIARULE aer_out_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_out_VIA7

VIARULE aer_in_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in_VIA4

VIARULE aer_in_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in_VIA3

VIARULE aer_in_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END aer_in_VIA2

VIARULE aer_in_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in_VIA1

VIARULE aer_in_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END aer_in_VIA0

VIARULE M3_M2$$219228204 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$219228204

VIARULE M3_M2$$193586220 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193586220

VIARULE M2_M1$$193575980 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193575980

VIARULE M2_M1$$193667116 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193667116

VIARULE M1_POLY1$$224275500 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$224275500

VIARULE M1_POLY1$$190326828 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$190326828

VIARULE M4_M3$$193802284 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M4_M3$$193802284

VIARULE M3_M2$$193580076 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2$$193580076

VIARULE M1_POLY1$$190324780 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.4 BY 0.4 ;
END M1_POLY1$$190324780

VIARULE M2_M1$$193805356 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1$$193805356

VIARULE M2_M1$$193668140 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193668140

VIARULE M2_M1$$212048940 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$212048940

VIARULE M2_M1$$193658924 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193658924

VIARULE M2_M1$$193808428 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193808428

VIARULE M2_M1$$193807404 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193807404

VIARULE M2_M1$$219750444 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$219750444

VIARULE M2_M1$$224472108 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$224472108

VIARULE M4_M3$$212047916 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$212047916

VIARULE M3_M2$$193581100 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193581100

VIARULE M3_M2$$224854060 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$224854060

VIARULE M2_M1$$193665068 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193665068

VIARULE M4_M3$$228254764 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$228254764

VIARULE M3_M2$$193587244 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193587244

VIARULE M4_M3$$224272428 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$224272428

VIARULE M2_M1$$193574956 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193574956

VIARULE M3_M2$$224471084 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$224471084

VIARULE M2_M1$$224841772 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$224841772

VIARULE M1_POLY1$$224473132 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$224473132

VIARULE M2_M1$$193660972 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193660972

VIARULE M2_M1$$224460844 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$224460844

VIARULE M1_POLY1$$224278572 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 1 ;
END M1_POLY1$$224278572

VIARULE M1_POLY1$$224848940 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 1 ;
END M1_POLY1$$224848940

VIARULE M2_M1$$193965100 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193965100

VIARULE M1_POLY1$$224191532 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M1_POLY1$$224191532

VIARULE M1_POLY1$$224190508 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$224190508

VIARULE M1_POLY1$$224189484 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$224189484

VIARULE M1_POLY1$$219225132 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$219225132

VIARULE M1_POLY1$$224188460 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$224188460

VIARULE M1_POLY1$$224277548 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$224277548

VIARULE M1_POLY1$$219741228 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 1 ;
END M1_POLY1$$219741228

VIARULE M1_POLY1$$224276524 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$224276524

VIARULE M1_POLY1$$190327852 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$190327852

VIARULE M3_M2$$241927212 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$241927212

VIARULE M4_M3$$222153772 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$222153772

VIARULE M3_M2$$193798188 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193798188

VIARULE M3_M2$$223323180 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$223323180

VIARULE M2_M1$$223320108 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$223320108

VIARULE M2_M1$$223319084 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$223319084

VIARULE M4_M3$$232261676 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$232261676

VIARULE M3_M2$$232412204 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$232412204

VIARULE M2_M1$$232411180 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232411180

VIARULE M2_M1$$193811500 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193811500

VIARULE M4_M3$$193957932 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 2 BY 1 ;
END M4_M3$$193957932

VIARULE M4_M3$$193956908 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 2 BY 1 ;
END M4_M3$$193956908

VIARULE M4_M3$$193955884 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 2 BY 1 ;
END M4_M3$$193955884

VIARULE M3_M2$$193954860 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 2 BY 1 ;
END M3_M2$$193954860

VIARULE M3_M2$$200606764 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 2 BY 1 ;
END M3_M2$$200606764

VIARULE M3_M2$$200605740 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 2 BY 1 ;
END M3_M2$$200605740

VIARULE M1_POLY1$$200604716 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 1 ;
END M1_POLY1$$200604716

VIARULE M2_M1$$200596524 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200596524

VIARULE M2_M1$$200593452 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200593452

VIARULE M2_M1$$193966124 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193966124

VIARULE M2_M1$$193964076 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193964076

VIARULE M2_M1$$193963052 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193963052

VIARULE M2_M1$$200598572 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200598572

VIARULE M1_POLY1$$193962028 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$193962028

VIARULE M2_M1$$200602668 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200602668

VIARULE M2_M1$$200601644 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200601644

VIARULE M2_M1$$200600620 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200600620

VIARULE M2_M1$$200599596 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200599596

VIARULE M1_POLY1$$200597548 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$200597548

VIARULE M3_M2$$229054508 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$229054508

VIARULE M2_M1$$193670188 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193670188

VIARULE M2_M1$$232266796 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232266796

VIARULE M2_M1$$232267820 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232267820

VIARULE M3_M2$$193583148 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193583148

VIARULE M3_M2$$232268844 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$232268844

VIARULE M3_M2$$232269868 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$232269868

VIARULE M4_M3$$232270892 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$232270892

VIARULE M4_M3$$232271916 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$232271916

VIARULE M4_M3$$231682092 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$231682092

VIARULE M2_M1$$232151084 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232151084

VIARULE M3_M2$$232276012 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$232276012

VIARULE M4_M3$$232272940 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$232272940

VIARULE M2_M1$$193657900 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193657900

VIARULE M3_M2$$228406316 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$228406316

VIARULE M3_M2$$232277036 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$232277036

VIARULE M2_M1$$231687212 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$231687212

VIARULE M2_M1$$231686188 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$231686188

VIARULE M2_M1$$231685164 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$231685164

VIARULE M3_M2$$229050412 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$229050412

VIARULE M1_POLY1$$227875884 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 1 ;
END M1_POLY1$$227875884

VIARULE M1_POLY1$$228018220 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$228018220

VIARULE M1_POLY1$$228019244 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 1 ;
END M1_POLY1$$228019244

VIARULE M1_POLY1$$233962540 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 1 ;
END M1_POLY1$$233962540

VIARULE M1_POLY1$$243994668 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 1 ;
END M1_POLY1$$243994668

VIARULE M1_POLY1$$302988332 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 0.8 ;
END M1_POLY1$$302988332

VIARULE M2_M1$$193572908 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193572908

VIARULE M2_M1$$193573932 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193573932

VIARULE M2_M1$$193577004 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193577004

VIARULE M2_M1$$193578028 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193578028

VIARULE M2_M1$$193656876 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193656876

VIARULE M2_M1$$193659948 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193659948

VIARULE M2_M1$$193661996 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193661996

VIARULE M2_M1$$193663020 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193663020

VIARULE M2_M1$$193664044 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193664044

VIARULE M2_M1$$193666092 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193666092

VIARULE M2_M1$$193669164 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193669164

VIARULE M2_M1$$193671212 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193671212

VIARULE M2_M1$$193672236 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193672236

VIARULE M2_M1$$193806380 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193806380

VIARULE M2_M1$$193809452 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193809452

VIARULE M2_M1$$193810476 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$193810476

VIARULE M2_M1$$200592428 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200592428

VIARULE M2_M1$$200603692 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$200603692

VIARULE M2_M1$$219223084 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$219223084

VIARULE M2_M1$$219224108 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$219224108

VIARULE M2_M1$$227868716 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$227868716

VIARULE M2_M1$$227878956 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$227878956

VIARULE M2_M1$$227882028 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$227882028

VIARULE M2_M1$$228403244 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$228403244

VIARULE M2_M1$$228404268 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$228404268

VIARULE M2_M1$$229048364 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 2 BY 1 ;
END M2_M1$$229048364

VIARULE M2_M1$$232612908 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232612908

VIARULE M2_M1$$232875052 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232875052

VIARULE M2_M1$$232876076 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232876076

VIARULE M2_M1$$232877100 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232877100

VIARULE M2_M1$$232878124 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232878124

VIARULE M2_M1$$232879148 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232879148

VIARULE M2_M1$$232880172 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232880172

VIARULE M2_M1$$232881196 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232881196

VIARULE M2_M1$$232882220 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232882220

VIARULE M2_M1$$232884268 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$232884268

VIARULE M2_M1$$233301036 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233301036

VIARULE M2_M1$$233792556 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233792556

VIARULE M2_M1$$233793580 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233793580

VIARULE M2_M1$$233794604 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233794604

VIARULE M2_M1$$233795628 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233795628

VIARULE M2_M1$$233796652 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233796652

VIARULE M2_M1$$233797676 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233797676

VIARULE M2_M1$$233901100 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233901100

VIARULE M2_M1$$233902124 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$233902124

VIARULE M2_M1$$235796524 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$235796524

VIARULE M2_M1$$235801644 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$235801644

VIARULE M2_M1$$236016684 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$236016684

VIARULE M2_M1$$236448812 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$236448812

VIARULE M2_M1$$236449836 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$236449836

VIARULE M2_M1$$241926188 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$241926188

VIARULE M2_M1$$242606124 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$242606124

VIARULE M2_M1$$242608172 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$242608172

VIARULE M2_M1$$242609196 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$242609196

VIARULE M2_M1$$242610220 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$242610220

VIARULE M2_M1$$304280620 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$304280620

VIARULE M2_M1$$426922028 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$426922028

VIARULE M2_M1$$426925100 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$426925100

VIARULE M2_M1$$426926124 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1$$426926124

VIARULE M2_M1_1219 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1219

VIARULE M2_M1_1287 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1287

VIARULE M2_M1_1299 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1299

VIARULE M2_M1_1396 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1396

VIARULE M2_M1_1483 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1483

VIARULE M2_M1_1527 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1527

VIARULE M2_M1_1722 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1722

VIARULE M2_M1_1753 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1753

VIARULE M2_M1_1842 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1842

VIARULE M2_M1_1872 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_1872

VIARULE M2_M1_216 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_216

VIARULE M2_M1_266 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_266

VIARULE M2_M1_29671 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_29671

VIARULE M2_M1_29711 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_29711

VIARULE M2_M1_29766 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_29766

VIARULE M2_M1_321 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_321

VIARULE M2_M1_361 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_361

VIARULE M2_M1_892 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M2_M1_892

VIARULE M3_M2$$193582124 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193582124

VIARULE M3_M2$$193584172 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193584172

VIARULE M3_M2$$193585196 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193585196

VIARULE M3_M2$$193969196 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$193969196

VIARULE M3_M2$$200591404 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$200591404

VIARULE M3_M2$$212049964 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$212049964

VIARULE M3_M2$$219229228 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$219229228

VIARULE M3_M2$$219230252 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$219230252

VIARULE M3_M2$$227874860 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$227874860

VIARULE M3_M2$$228405292 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$228405292

VIARULE M3_M2$$233197612 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233197612

VIARULE M3_M2$$233198636 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233198636

VIARULE M3_M2$$233199660 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233199660

VIARULE M3_M2$$233200684 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233200684

VIARULE M3_M2$$233201708 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233201708

VIARULE M3_M2$$233202732 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233202732

VIARULE M3_M2$$233203756 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233203756

VIARULE M3_M2$$233204780 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233204780

VIARULE M3_M2$$233205804 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233205804

VIARULE M3_M2$$233206828 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233206828

VIARULE M3_M2$$233295916 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233295916

VIARULE M3_M2$$233296940 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233296940

VIARULE M3_M2$$233297964 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233297964

VIARULE M3_M2$$233298988 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233298988

VIARULE M3_M2$$233300012 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233300012

VIARULE M3_M2$$233798700 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233798700

VIARULE M3_M2$$233799724 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233799724

VIARULE M3_M2$$233800748 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233800748

VIARULE M3_M2$$233801772 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233801772

VIARULE M3_M2$$233802796 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233802796

VIARULE M3_M2$$233803820 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233803820

VIARULE M3_M2$$233804844 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233804844

VIARULE M3_M2$$233805868 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233805868

VIARULE M3_M2$$233806892 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233806892

VIARULE M3_M2$$233807916 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$233807916

VIARULE M3_M2$$236002348 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236002348

VIARULE M3_M2$$236003372 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236003372

VIARULE M3_M2$$236004396 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236004396

VIARULE M3_M2$$236017708 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236017708

VIARULE M3_M2$$236066860 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236066860

VIARULE M3_M2$$236442668 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236442668

VIARULE M3_M2$$236443692 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236443692

VIARULE M3_M2$$236444716 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236444716

VIARULE M3_M2$$236445740 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236445740

VIARULE M3_M2$$236446764 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236446764

VIARULE M3_M2$$236447788 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$236447788

VIARULE M3_M2$$241933356 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$241933356

VIARULE M3_M2$$302991404 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$302991404

VIARULE M3_M2$$426924076 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2$$426924076

VIARULE M3_M2_1218 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1218

VIARULE M3_M2_1286 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1286

VIARULE M3_M2_1300 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1300

VIARULE M3_M2_1395 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1395

VIARULE M3_M2_1484 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1484

VIARULE M3_M2_1528 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1528

VIARULE M3_M2_1723 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1723

VIARULE M3_M2_1754 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1754

VIARULE M3_M2_1841 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1841

VIARULE M3_M2_1871 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_1871

VIARULE M3_M2_215 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_215

VIARULE M3_M2_265 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_265

VIARULE M3_M2_29672 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_29672

VIARULE M3_M2_29710 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_29710

VIARULE M3_M2_29767 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_29767

VIARULE M3_M2_322 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_322

VIARULE M3_M2_362 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_362

VIARULE M3_M2_891 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END M3_M2_891

VIARULE M4_M3$$193799212 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$193799212

VIARULE M4_M3$$193803308 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$193803308

VIARULE M4_M3$$229053484 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$229053484

VIARULE M4_M3$$233207852 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233207852

VIARULE M4_M3$$233208876 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233208876

VIARULE M4_M3$$233209900 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233209900

VIARULE M4_M3$$233210924 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233210924

VIARULE M4_M3$$233886764 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233886764

VIARULE M4_M3$$233887788 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233887788

VIARULE M4_M3$$233888812 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233888812

VIARULE M4_M3$$233889836 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233889836

VIARULE M4_M3$$233890860 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233890860

VIARULE M4_M3$$233891884 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233891884

VIARULE M4_M3$$233892908 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233892908

VIARULE M4_M3$$233893932 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233893932

VIARULE M4_M3$$233894956 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233894956

VIARULE M4_M3$$233895980 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233895980

VIARULE M4_M3$$233897004 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233897004

VIARULE M4_M3$$233898028 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233898028

VIARULE M4_M3$$233899052 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233899052

VIARULE M4_M3$$233900076 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233900076

VIARULE M4_M3$$233958444 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233958444

VIARULE M4_M3$$233963564 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233963564

VIARULE M4_M3$$233964588 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233964588

VIARULE M4_M3$$233965612 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233965612

VIARULE M4_M3$$233966636 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233966636

VIARULE M4_M3$$233967660 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233967660

VIARULE M4_M3$$233968684 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233968684

VIARULE M4_M3$$233969708 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233969708

VIARULE M4_M3$$233970732 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$233970732

VIARULE M4_M3$$235795500 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$235795500

VIARULE M4_M3$$235799596 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$235799596

VIARULE M4_M3$$235800620 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$235800620

VIARULE M4_M3$$235802668 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$235802668

VIARULE M4_M3$$235803692 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$235803692

VIARULE M4_M3$$236005420 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236005420

VIARULE M4_M3$$236006444 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236006444

VIARULE M4_M3$$236007468 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236007468

VIARULE M4_M3$$236008492 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236008492

VIARULE M4_M3$$236009516 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236009516

VIARULE M4_M3$$236010540 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236010540

VIARULE M4_M3$$236011564 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236011564

VIARULE M4_M3$$236012588 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236012588

VIARULE M4_M3$$236013612 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236013612

VIARULE M4_M3$$236014636 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236014636

VIARULE M4_M3$$236015660 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236015660

VIARULE M4_M3$$236064812 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236064812

VIARULE M4_M3$$236065836 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236065836

VIARULE M4_M3$$236067884 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236067884

VIARULE M4_M3$$236068908 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236068908

VIARULE M4_M3$$236080172 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236080172

VIARULE M4_M3$$236450860 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236450860

VIARULE M4_M3$$236451884 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236451884

VIARULE M4_M3$$236452908 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236452908

VIARULE M4_M3$$236453932 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236453932

VIARULE M4_M3$$236454956 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236454956

VIARULE M4_M3$$236455980 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236455980

VIARULE M4_M3$$236541996 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236541996

VIARULE M4_M3$$236543020 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$236543020

VIARULE M4_M3$$242607148 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$242607148

VIARULE M4_M3$$243494956 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$243494956

VIARULE M4_M3$$243507244 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$243507244

VIARULE M4_M3$$391955500 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$391955500

VIARULE M4_M3$$391956524 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$391956524

VIARULE M4_M3$$426923052 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL4 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3$$426923052

VIARULE prog_periph_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END prog_periph_VIA7

VIARULE prog_periph_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END prog_periph_VIA6

VIARULE prog_periph_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END prog_periph_VIA5

VIARULE prog_periph_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END prog_periph_VIA4

VIARULE prog_periph_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END prog_periph_VIA3

VIARULE prog_periph_VIA2 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END prog_periph_VIA2

VIARULE prog_periph_VIA1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END prog_periph_VIA1

VIARULE prog_periph_VIA0 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.5 BY 0.5 ;
END prog_periph_VIA0

VIARULE openMSP430_VIA7 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.175 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.175 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 0.95 ;
END openMSP430_VIA7

VIARULE openMSP430_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END openMSP430_VIA6

VIARULE openMSP430_VIA5 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.175 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.175 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 0.95 ;
END openMSP430_VIA5

VIARULE openMSP430_VIA4 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.375 ;
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.375 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 0.95 ;
END openMSP430_VIA4

VIARULE openMSP430_VIA3 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER METAL2 ;
    ENCLOSURE 0.375 0.625 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END openMSP430_VIA3

VIARULE dacbank_periph_VIA6 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER METAL2 ;
    ENCLOSURE 0.35 0.425 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 0.95 BY 0.95 ;
END dacbank_periph_VIA6

