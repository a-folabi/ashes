module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(6), .GND_b_1_row_4(net1606[0:6]), .Vs_b_0_row_4(net112[0:6]), .Vs_b_1_row_4(net113[0:6]), .VINJ_b_1_row_4(net1612[0:6]), .Vsel_b_0_row_4(net1576[0:6]), .Vsel_b_1_row_4(net1577[0:6]), .Vg_b_0_row_4(net1588[0:6]), .Vg_b_1_row_4(net1589[0:6]), .VTUN_brow_4(net1600[0:6]), .Vd_Rl_0_col_0(net1941[0:5]), .Vd_Rl_1_col_0(net1942[0:5]), .Vd_Rl_2_col_0(net1943[0:5]), .Vd_Rl_3_col_0(net1944[0:5]), .Vd_Pl_0_col_0(net1772[0:5]), .Vd_Pl_1_col_0(net1773[0:5]), .Vd_Pl_2_col_0(net1774[0:5]), .Vd_Pl_3_col_0(net1775[0:5]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(6), .GND_b_1_row_4(net1645[0:6]), .Vs_b_0_row_4(net237[0:6]), .Vs_b_1_row_4(net236[0:6]), .VINJ_b_1_row_4(net1644[0:6]), .Vsel_b_0_row_4(net1646[0:6]), .Vsel_b_1_row_4(net1648[0:6]), .Vg_b_0_row_4(net1647[0:6]), .Vg_b_1_row_4(net1649[0:6]), .VTUN_brow_4(net1643[0:6]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(22), .matrix_row(5), .matrix_col(1), .A_0_col_0(net1975[0:5]), .A_1_col_0(net1976[0:5]), .A_2_col_0(net1977[0:5]), .A_3_col_0(net1978[0:5]), .Prog_brow_4(net1934[0:1]), .VDD_brow_4(net1913[0:1]), .GND_brow_4(net1645[5:6]), .Progrow_0(net1934[0:1]));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(6), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1622[0:1]), .Vsel_b_0_row_4(net1625[0:1]), .Vsel_b_1_row_4(net1626[0:1]), .Vg_b_0_row_4(net1627[0:1]), .Vg_b_1_row_4(net1628[0:1]), .VTUN_brow_4(net1623[0:1]), .GND_b_1_row_4(net1624[0:1]));
	S_BLOCK_BUFFER I__4 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__5 (.island_num(0), .row(0), .col(8), .matrix_row(4), .matrix_col(1), .n_0_row_0(net1882[0:1]), .n_1_row_0(net1883[0:1]), .n_2_row_0(net1884[0:1]), .n_3_row_0(net1885[0:1]));
	S_BLOCK_CONN_PINS I__6 (.island_num(0), .row(4), .col(8), .matrix_row(1), .matrix_col(1), .s_0_row_0(net1914), .s_1_row_0(net1915), .s_2_row_0(net1916), .s_3_row_0(net1917));
	S_BLOCK_SPACE_UP_PINS I__7 (.island_num(0), .row(0), .col(9), .matrix_row(3), .matrix_col(1), .n_0_row_0(net1886[0:1]), .n_1_row_0(net1887[0:1]), .n_2_row_0(net1888[0:1]), .n_3_row_0(net1889[0:1]));
	S_BLOCK_CONN_PINS I__8 (.island_num(0), .row(3), .col(9), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__9 (.island_num(0), .row(4), .col(9), .matrix_row(1), .matrix_col(1), .s_0_row_0(net1918), .s_1_row_0(net1919), .s_2_row_0(net1920), .s_3_row_0(net1921));
	S_BLOCK_SPACE_UP_PINS I__10 (.island_num(0), .row(0), .col(10), .matrix_row(2), .matrix_col(1), .n_0_row_0(net1890[0:1]), .n_1_row_0(net1891[0:1]), .n_2_row_0(net1892[0:1]), .n_3_row_0(net1893[0:1]));
	S_BLOCK_CONN_PINS I__11 (.island_num(0), .row(2), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__12 (.island_num(0), .row(3), .col(10), .matrix_row(2), .matrix_col(1), .s_0_row_1(net1922[0:1]), .s_1_row_1(net1923[0:1]), .s_2_row_1(net1924[0:1]), .s_3_row_1(net1925[0:1]));
	S_BLOCK_SPACE_UP_PINS I__13 (.island_num(0), .row(0), .col(11), .matrix_row(1), .matrix_col(1), .n_0_row_0(net1894), .n_1_row_0(net1895), .n_2_row_0(net1896), .n_3_row_0(net1897));
	S_BLOCK_CONN_PINS I__14 (.island_num(0), .row(1), .col(11), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__15 (.island_num(0), .row(2), .col(11), .matrix_row(3), .matrix_col(1), .s_0_row_2(net1926[0:1]), .s_1_row_2(net1927[0:1]), .s_2_row_2(net1928[0:1]), .s_3_row_2(net1929[0:1]));
	S_BLOCK_CONN_PINS I__16 (.island_num(0), .row(0), .col(12), .matrix_row(1), .matrix_col(1), .n_0_row_0(net1898), .n_1_row_0(net1899), .n_2_row_0(net1900), .n_3_row_0(net1901));
	S_BLOCK_SPACE_DOWN_PINS I__17 (.island_num(0), .row(1), .col(12), .matrix_row(4), .matrix_col(1), .s_0_row_3(net1930[0:1]), .s_1_row_3(net1931[0:1]), .s_2_row_3(net1932[0:1]), .s_3_row_3(net1933[0:1]));
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(13), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1629[0:1]), .Vsel_b_0_row_4(net1632[0:1]), .Vsel_b_1_row_4(net1633[0:1]), .Vg_b_0_row_4(net1634[0:1]), .Vg_b_1_row_4(net1635[0:1]), .VTUN_brow_4(net1630[0:1]), .GND_b_1_row_4(net1631[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net1636[0:1]), .Vsel_b_0_row_4(net1639[0:1]), .Vsel_b_1_row_4(net1640[0:1]), .Vg_b_0_row_4(net1641[0:1]), .Vg_b_1_row_4(net1642[0:1]), .VTUN_brow_4(net1637[0:1]), .GND_b_1_row_4(net1638[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(5), .decode_n1_VGRUN_2_(net1878[0]), .decode_n1_VGRUN_3_(net1879[0]), .decode_n2_VGRUN_0_(net1880[0]), .decode_n2_VGRUN_1_(net1881[0]), .decode_n5_VGRUN_2_(net1961[0]), .decode_n5_VGRUN_3_(net1962[0]), .decode_n6_VGRUN_0_(net1963[0]), .decode_n6_VGRUN_1_(net1964[0]), .decode_n4_n0_RUN_OUT_0_(net1748[0]), .decode_n4_n0_RUN_OUT_1_(net1749[0]), .decode_n4_n0_RUN_OUT_2_(net1750[0]), .decode_n4_n0_RUN_OUT_3_(net1751[0]), .decode_n4_n1_RUN_OUT_0_(net1752[0]), .decode_n4_n1_RUN_OUT_1_(net1753[0]), .decode_n4_n1_RUN_OUT_2_(net1740), .decode_n4_n1_RUN_OUT_3_(net1741), .decode_n4_n2_RUN_OUT_0_(net1742), .decode_n4_n2_RUN_OUT_1_(net1743), .decode_n4_n2_RUN_OUT_2_(net1754[0]), .decode_n4_n2_RUN_OUT_3_(net1755[0]), .decode_n4_n3_RUN_OUT_0_(net1756[0]), .decode_n4_n3_RUN_OUT_1_(net1757[0]), .decode_n4_n3_RUN_OUT_2_(net1758[0]), .decode_n4_n3_RUN_OUT_3_(net1759[0]), .decode_n4_n4_RUN_OUT_0_(net1760[0]), .decode_n4_n4_RUN_OUT_1_(net1761[0]), .decode_n4_n4_RUN_OUT_2_(net1762[0]), .decode_n4_n4_RUN_OUT_3_(net1763[0]), .decode_n4_n5_RUN_OUT_0_(net1764[0]), .decode_n4_n5_RUN_OUT_1_(net1765[0]), .decode_n4_n5_RUN_OUT_2_(net1744), .decode_n4_n5_RUN_OUT_3_(net1745), .decode_n4_n6_RUN_OUT_0_(net1746), .decode_n4_n6_RUN_OUT_1_(net1747), .decode_n4_n6_RUN_OUT_2_(net1766[0]), .decode_n4_n6_RUN_OUT_3_(net1767[0]), .decode_n4_n7_RUN_OUT_0_(net1768[0]), .decode_n4_n7_RUN_OUT_1_(net1769[0]), .decode_n4_n7_RUN_OUT_2_(net1770[0]), .decode_n4_n7_RUN_OUT_3_(net1771[0]), .decode_n4_n0_OUT_0_(net1686), .decode_n4_n0_OUT_1_(net1687), .decode_n4_n0_OUT_2_(net1690), .decode_n4_n0_OUT_3_(net1691), .decode_n4_n1_OUT_0_(net1694), .decode_n4_n1_OUT_1_(net1695), .decode_n4_n1_OUT_2_(net1698), .decode_n4_n1_OUT_3_(net1699), .decode_n4_n2_OUT_0_(net1702), .decode_n4_n2_OUT_1_(net1703), .decode_n4_n2_OUT_2_(net1706), .decode_n4_n2_OUT_3_(net1707), .decode_n4_n3_OUT_0_(net1710), .decode_n4_n3_OUT_1_(net1711), .decode_n4_n4_OUT_0_(net1714), .decode_n4_n4_OUT_1_(net1715), .decode_n4_n4_OUT_2_(net1718), .decode_n4_n4_OUT_3_(net1719), .decode_n4_n5_OUT_0_(net1722), .decode_n4_n5_OUT_1_(net1723), .decode_n4_n5_OUT_2_(net1726), .decode_n4_n5_OUT_3_(net1727), .decode_n4_n6_OUT_0_(net1730), .decode_n4_n6_OUT_1_(net1731), .decode_n4_n6_OUT_2_(net1734), .decode_n4_n6_OUT_3_(net1735), .decode_n4_n7_OUT_0_(net1738), .decode_n4_n7_OUT_1_(net1739), .decode_n0_ENABLE(net1902), .decode_n4_n0_VINJ_b_0_(net1684), .decode_n4_n0_VINJ_b_1_(net1688), .decode_n4_n1_VINJ_b_0_(net1692), .decode_n4_n1_VINJ_b_1_(net1696), .decode_n4_n2_VINJ_b_0_(net1700), .decode_n4_n2_VINJ_b_1_(net1704), .decode_n4_n3_VINJ_b_0_(net1708), .decode_n4_n4_VINJ_b_0_(net1712), .decode_n4_n4_VINJ_b_1_(net1716), .decode_n4_n5_VINJ_b_0_(net1720), .decode_n4_n5_VINJ_b_1_(net1724), .decode_n4_n6_VINJ_b_0_(net1728), .decode_n4_n6_VINJ_b_1_(net1732), .decode_n4_n7_VINJ_b_0_(net1736), .decode_n4_n0_GND_b_0_(net1685), .decode_n4_n0_GND_b_1_(net1689), .decode_n4_n1_GND_b_0_(net1693), .decode_n4_n1_GND_b_1_(net1697), .decode_n4_n2_GND_b_0_(net1701), .decode_n4_n2_GND_b_1_(net1705), .decode_n4_n3_GND_b_0_(net1709), .decode_n4_n4_GND_b_0_(net1713), .decode_n4_n4_GND_b_1_(net1717), .decode_n4_n5_GND_b_0_(net1721), .decode_n4_n5_GND_b_1_(net1725), .decode_n4_n6_GND_b_0_(net1729), .decode_n4_n6_GND_b_1_(net1733), .decode_n4_n7_GND_b_0_(net1737), .decode_n0_VINJV(net1909), .decode_n0_GNDV(net1911));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(22), .switch_n3_VPWR_0_(net1740), .switch_n3_VPWR_1_(net1741), .switch_n4_VPWR_0_(net1742), .switch_n4_VPWR_1_(net1743), .switch_n17_VPWR_0_(net1744), .switch_n17_VPWR_1_(net1745), .switch_n18_VPWR_0_(net1746), .switch_n18_VPWR_1_(net1747), .switch_n0_RUN_IN_0_(net1877), .switch_n0_RUN_IN_1_(net1877), .switch_n1_RUN_IN_0_(net1877), .switch_n1_RUN_IN_1_(net1877), .switch_n2_RUN_IN_0_(net1877), .switch_n2_RUN_IN_1_(net1877), .switch_n3_RUN_IN_0_(net1877), .switch_n3_RUN_IN_1_(net1877), .switch_n4_RUN_IN_0_(net1877), .switch_n4_RUN_IN_1_(net1877), .switch_n5_RUN_IN_0_(net1877), .switch_n5_RUN_IN_1_(net1877), .switch_n6_RUN_IN_0_(net1877), .switch_n6_RUN_IN_1_(net1877), .switch_n13_RUN_IN_0_(net1877), .switch_n13_RUN_IN_1_(net1877), .switch_n15_RUN_IN_0_(net1877), .switch_n15_RUN_IN_1_(net1877), .switch_n16_RUN_IN_0_(net1877), .switch_n16_RUN_IN_1_(net1877), .switch_n17_RUN_IN_0_(net1877), .switch_n17_RUN_IN_1_(net1877), .switch_n18_RUN_IN_0_(net1877), .switch_n18_RUN_IN_1_(net1877), .switch_n19_RUN_IN_0_(net1877), .switch_n19_RUN_IN_1_(net1877), .switch_n20_RUN_IN_0_(net1877), .switch_n20_RUN_IN_1_(net1877), .switch_n21_RUN_IN_0_(net1877), .switch_n21_RUN_IN_1_(net1877), .switch_n0_GND_T(net1685), .switch_n1_GND_T(net1689), .switch_n2_GND_T(net1693), .switch_n3_GND_T(net1697), .switch_n4_GND_T(net1701), .switch_n5_GND_T(net1705), .switch_n6_GND_T(net1709), .switch_n14_GND_T(net1713), .switch_n15_GND_T(net1717), .switch_n16_GND_T(net1721), .switch_n17_GND_T(net1725), .switch_n18_GND_T(net1729), .switch_n19_GND_T(net1733), .switch_n20_GND_T(net1737), .switch_n0_VTUN_T(net1966[0]), .switch_n0_decode_0_(net1686), .switch_n0_decode_1_(net1687), .switch_n1_decode_0_(net1690), .switch_n1_decode_1_(net1691), .switch_n2_decode_0_(net1694), .switch_n2_decode_1_(net1695), .switch_n3_decode_0_(net1698), .switch_n3_decode_1_(net1699), .switch_n4_decode_0_(net1702), .switch_n4_decode_1_(net1703), .switch_n5_decode_0_(net1706), .switch_n5_decode_1_(net1707), .switch_n6_decode_0_(net1710), .switch_n6_decode_1_(net1711), .switch_n14_decode_0_(net1714), .switch_n14_decode_1_(net1715), .switch_n15_decode_0_(net1718), .switch_n15_decode_1_(net1719), .switch_n16_decode_0_(net1722), .switch_n16_decode_1_(net1723), .switch_n17_decode_0_(net1726), .switch_n17_decode_1_(net1727), .switch_n18_decode_0_(net1730), .switch_n18_decode_1_(net1731), .switch_n19_decode_0_(net1734), .switch_n19_decode_1_(net1735), .switch_n20_decode_0_(net1738), .switch_n20_decode_1_(net1739), .switch_n0_VINJ_T(net1684), .switch_n1_VINJ_T(net1688), .switch_n2_VINJ_T(net1692), .switch_n3_VINJ_T(net1696), .switch_n4_VINJ_T(net1700), .switch_n5_VINJ_T(net1704), .switch_n6_VINJ_T(net1708), .switch_n14_VINJ_T(net1712), .switch_n15_VINJ_T(net1716), .switch_n16_VINJ_T(net1720), .switch_n17_VINJ_T(net1724), .switch_n18_VINJ_T(net1728), .switch_n19_VINJ_T(net1732), .switch_n20_VINJ_T(net1736), .switch_n0_RUN(net1935), .switch_n0_vgsel_r(net1936));
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5), .decode_n0_IN_0_(net1974), .decode_n0_IN_1_(net1973), .decode_n0_IN_2_(net1972), .decode_n0_IN_3_(net1971), .decode_n0_IN_4_(net1970), .decode_n0_ENABLE(net2000));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select), .switch_n0_prog_drainrail(net1903), .switch_n0_run_drainrail(net1904), .switch_n0_VINJ(net1910), .switch_n0_GND(net1912));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch), .switch_n0_PR_0_(net1772[0]), .switch_n0_PR_1_(net1773[0]), .switch_n0_PR_2_(net1774[0]), .switch_n0_PR_3_(net1775[0]), .switch_n1_PR_0_(net1772[1]), .switch_n1_PR_1_(net1773[1]), .switch_n1_PR_2_(net1774[1]), .switch_n1_PR_3_(net1775[1]), .switch_n2_PR_0_(net1772[2]), .switch_n2_PR_1_(net1773[2]), .switch_n2_PR_2_(net1774[2]), .switch_n2_PR_3_(net1775[2]), .switch_n3_PR_0_(net1772[3]), .switch_n3_PR_1_(net1773[3]), .switch_n3_PR_2_(net1774[3]), .switch_n3_PR_3_(net1775[3]), .switch_n4_PR_0_(net1772[4]), .switch_n4_PR_1_(net1773[4]), .switch_n4_PR_2_(net1774[4]), .switch_n4_PR_3_(net1775[4]), .switch_n0_In_0_(net1941[0]), .switch_n0_In_1_(net1942[0]), .switch_n0_In_2_(net1943[0]), .switch_n0_In_3_(net1944[0]), .switch_n1_In_0_(net1941[1]), .switch_n1_In_1_(net1942[1]), .switch_n1_In_2_(net1943[1]), .switch_n1_In_3_(net1944[1]), .switch_n2_In_0_(net1941[2]), .switch_n2_In_1_(net1942[2]), .switch_n2_In_2_(net1943[2]), .switch_n2_In_3_(net1944[2]), .switch_n3_In_0_(net1941[3]), .switch_n3_In_1_(net1942[3]), .switch_n3_In_2_(net1943[3]), .switch_n3_In_3_(net1944[3]), .switch_n4_In_0_(net1941[4]), .switch_n4_In_1_(net1942[4]), .switch_n4_In_2_(net1943[4]), .switch_n4_In_3_(net1944[4]), .switch_n0_VDD(net1910), .switch_n0_GND(net1912), .switch_n0_RUN(net1935));
	none switch_ind(.island_num(0), .direction(horizontal), .col(7));
	none switch_ind(.island_num(0), .direction(horizontal), .col(8));
	none switch_ind(.island_num(0), .direction(horizontal), .col(9));
	none switch_ind(.island_num(0), .direction(horizontal), .col(10));
	none switch_ind(.island_num(0), .direction(horizontal), .col(11));
	none switch_ind(.island_num(0), .direction(horizontal), .col(12));
	none switch_ind(.island_num(0), .direction(horizontal), .col(14));


	/* Island 1 */
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__0 (.island_num(1), .row(0), .col(0), .matrix_row(1), .matrix_col(8));
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(5), .matrix_col(8), .GND_b_0_row_4(net893[0:8]), .GND_b_1_row_4(net894[0:8]), .Vs_b_0_row_4(net903[0:8]), .Vs_b_1_row_4(net904[0:8]), .VINJ_b_0_row_4(net907[0:8]), .VINJ_b_1_row_4(net908[0:8]), .Vsel_b_0_row_4(net911[0:8]), .Vsel_b_1_row_4(net912[0:8]), .Vg_b_0_row_4(net915[0:8]), .Vg_b_1_row_4(net916[0:8]), .VTUN_brow_4(net919[0:8]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(8), .matrix_row(1), .matrix_col(6));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(8), .matrix_row(4), .matrix_col(6));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(5), .col(8), .matrix_row(1), .matrix_col(6));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(14), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1523), .P_1_row_0(net1524), .A_0_row_0(net1525), .A_1_row_0(net1526), .A_2_row_0(net1527), .A_3_row_0(net1528), .Progrow_0(net1873), .VDDrow_0(net1913[0]), .GNDrow_0(net1645[5]));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(14), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1536), .P_1_row_0(net1537), .A_0_row_0(net1538), .A_1_row_0(net1539), .A_2_row_0(net1540), .A_3_row_0(net1541));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(14), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1550), .A_1_row_0(net1551), .A_2_row_0(net1552), .A_3_row_0(net1553));
	TSMC350nm_4TGate_ST_BMatrix I__8 (.island_num(1), .row(3), .col(14), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1559), .A_1_row_0(net1560), .A_2_row_0(net1561), .A_3_row_0(net1562));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(14), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1568), .A_1_row_0(net1569), .A_2_row_0(net1570), .A_3_row_0(net1571));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(14), .matrix_row(1), .matrix_col(1), .Prog_brow_0(net1876[0]), .VDD_brow_0(net1875[0]), .GND_brow_0(net1874[0]));
	TSMC350nm_OutMtrx_IndrctSwcs I__11 (.island_num(1), .row(7), .col(8), .matrix_row(1), .matrix_col(6));
	TSMC350nm_4x2_Indirect I__12 (.island_num(1), .row(8), .col(8), .matrix_row(2), .matrix_col(6), .Vd_Rl_0_col_0(net1387[0:2]), .Vd_Rl_1_col_0(net1388[0:2]), .Vd_Rl_2_col_0(net1389[0:2]), .Vd_Rl_3_col_0(net1390[0:2]), .Vd_Pl_0_col_0(net1391[0:2]), .Vd_Pl_1_col_0(net1392[0:2]), .Vd_Pl_2_col_0(net1393[0:2]), .Vd_Pl_3_col_0(net1394[0:2]));
	TSMC350nm_4TGate_ST_BMatrix I__13 (.island_num(1), .row(8), .col(14), .matrix_row(2), .matrix_col(1), .A_0_col_0(net1905[0:2]), .A_1_col_0(net1906[0:2]), .A_2_col_0(net1907[0:2]), .A_3_col_0(net1908[0:2]), .Progrow_0(net1876[0:1]), .VDDrow_0(net1875[0:1]), .GNDrow_0(net1874[0:1]));
	TSMC350nm_TA2Cell_NoFG cab_device_14 (.island_num(1), .row(2), .col(15), .VD_P_0_(net1523), .VD_P_1_(net1524), .VIN1_PLUS(net1525), .VIN1_MINUS(net1526), .VIN2_PLUS(net1527), .VIN2_MINUS(net1528), .OUTPUT_0_(net1529[0]), .OUTPUT_1_(net1530[0]), .VTUN(net1531), .Vg(net1532), .Vsel(net1533), .VINJ(net1534), .GND(net1535), .VPWR(net1969[0]), .VTUN_b(net1544), .Vg_b(net1545), .Vsel_b(net1546), .VINJ_b(net1547), .GND_b(net1548), .VPWR_b(net1549));
	TSMC350nm_TA2Cell_NoFG cab_device_15 (.island_num(1), .row(3), .col(15), .VD_P_0_(net1536), .VD_P_1_(net1537), .VIN1_PLUS(net1538), .VIN1_MINUS(net1539), .VIN2_PLUS(net1540), .VIN2_MINUS(net1541), .OUTPUT_0_(net1542[0]), .OUTPUT_1_(net1543[0]), .VTUN(net1544), .Vg(net1545), .Vsel(net1546), .VINJ(net1547), .GND(net1548), .VPWR(net1549), .GND_b(net1558), .VPWR_b(net1557));
	TSMC350nm_TGate_2nMirror cab_device_16 (.island_num(1), .row(4), .col(15), .IN_CM_0_(net1550), .IN_CM_1_(net1551), .SelN(net1552), .IN_TG(net1553), .OUT_CM_0_(net1554[0]), .OUT_CM_1_(net1555[0]), .OUT_TG(net1556[0]), .VPWR(net1557), .GND(net1558), .VPWR_b(net1566), .GND_b(net1567));
	TSMC350nm_TGate_2nMirror cab_device_17 (.island_num(1), .row(5), .col(15), .IN_CM_0_(net1559), .IN_CM_1_(net1560), .SelN(net1561), .IN_TG(net1562), .OUT_CM_0_(net1563[0]), .OUT_CM_1_(net1564[0]), .OUT_TG(net1565[0]), .VPWR(net1566), .GND(net1567), .VPWR_b(net1574), .GND_b(net1575));
	TSMC350nm_NandPfets cab_device_18 (.island_num(1), .row(6), .col(15), .GATE_N(net1568), .SOURCE_N(net1569), .GATE_P(net1570), .SOURCE_P(net1571), .DRAIN_N(net1572[0]), .DRAIN_P(net1573[0]), .VPWR(net1574), .GND(net1575));
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6), .decode_n0_IN_0_(net1999), .decode_n0_IN_1_(net1998), .decode_n0_IN_2_(net1997), .decode_n0_IN_3_(net1996), .decode_n0_IN_4_(net1995), .decode_n0_ENABLE(net2000));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(1), .direction(vertical), .num(10), .type(drain_select), .switch_n0_prog_drainrail(net1903), .switch_n0_run_drainrail(net1904));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(10), .type(prog_switch), .switch_n6_PR_0_(net1857[0]), .switch_n6_PR_1_(net1861[0]), .switch_n6_PR_2_(net1865[0]), .switch_n6_PR_3_(net1869[0]), .switch_n6_In_0_(net1856[0]), .switch_n6_In_1_(net1860[0]), .switch_n6_In_2_(net1864[0]), .switch_n6_In_3_(net1868[0]), .switch_n0_RUN(net1935));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(16), .switch_n0_Input_0_(net1913[0]), .switch_n0_Input_1_(net1606[0]), .switch_n1_Input_0_(net112[1]), .switch_n1_Input_1_(net113[1]), .switch_n2_Input_0_(net112[2]), .switch_n2_Input_1_(net113[2]), .switch_n3_Input_0_(net237[0]), .switch_n7_Input_1_(net1855[0]), .switch_n8_Input_0_(net1529[0]), .switch_n8_Input_1_(net1530[0]), .switch_n9_Input_0_(net1542[0]), .switch_n9_Input_1_(net1543[0]), .switch_n10_Input_0_(net1554[0]), .switch_n10_Input_1_(net1555[0]), .switch_n11_Input_0_(net1556[0]), .switch_n11_Input_1_(net1563[0]), .switch_n12_Input_0_(net1564[0]), .switch_n12_Input_1_(net1565[0]), .switch_n13_Input_0_(net1572[0]), .switch_n13_Input_1_(net1573[0]), .switch_n0_GND(net1606[0]), .switch_n1_GND(net1606[1]), .switch_n2_GND(net1606[2]), .switch_n3_GND(net1606[3]), .switch_n4_GND(net1606[4]), .switch_n5_GND(net1606[5]), .switch_n6_GND(net1624[0]), .switch_n7_GND(net1631[0]), .switch_n8_GND(net1638[0]), .switch_n9_GND(net1645[0]), .switch_n10_GND(net1645[1]), .switch_n11_GND(net1645[2]), .switch_n12_GND(net1645[3]), .switch_n13_GND(net1645[4]), .switch_n14_GND(net1645[5]), .switch_n0_Vsel_0_(net1576[0]), .switch_n0_Vsel_1_(net1577[0]), .switch_n1_Vsel_0_(net1576[1]), .switch_n1_Vsel_1_(net1577[1]), .switch_n2_Vsel_0_(net1576[2]), .switch_n2_Vsel_1_(net1577[2]), .switch_n3_Vsel_0_(net1576[3]), .switch_n3_Vsel_1_(net1577[3]), .switch_n4_Vsel_0_(net1576[4]), .switch_n4_Vsel_1_(net1577[4]), .switch_n5_Vsel_0_(net1576[5]), .switch_n5_Vsel_1_(net1577[5]), .switch_n6_Vsel_0_(net1626[0]), .switch_n6_Vsel_1_(net1625[0]), .switch_n7_Vsel_0_(net1633[0]), .switch_n7_Vsel_1_(net1632[0]), .switch_n8_Vsel_0_(net1640[0]), .switch_n8_Vsel_1_(net1639[0]), .switch_n9_Vsel_0_(net1646[0]), .switch_n9_Vsel_1_(net1648[0]), .switch_n10_Vsel_0_(net1646[1]), .switch_n10_Vsel_1_(net1648[1]), .switch_n11_Vsel_0_(net1646[2]), .switch_n11_Vsel_1_(net1648[2]), .switch_n12_Vsel_0_(net1646[3]), .switch_n12_Vsel_1_(net1648[3]), .switch_n13_Vsel_0_(net1646[4]), .switch_n13_Vsel_1_(net1648[4]), .switch_n14_Vsel_0_(net1646[5]), .switch_n14_Vsel_1_(net1648[5]), .switch_n0_Vg_global_0_(net1588[0]), .switch_n0_Vg_global_1_(net1589[0]), .switch_n1_Vg_global_0_(net1588[1]), .switch_n1_Vg_global_1_(net1589[1]), .switch_n2_Vg_global_0_(net1588[2]), .switch_n2_Vg_global_1_(net1589[2]), .switch_n3_Vg_global_0_(net1588[3]), .switch_n3_Vg_global_1_(net1589[3]), .switch_n4_Vg_global_0_(net1588[4]), .switch_n4_Vg_global_1_(net1589[4]), .switch_n5_Vg_global_0_(net1588[5]), .switch_n5_Vg_global_1_(net1589[5]), .switch_n6_Vg_global_0_(net1628[0]), .switch_n6_Vg_global_1_(net1627[0]), .switch_n7_Vg_global_0_(net1635[0]), .switch_n7_Vg_global_1_(net1634[0]), .switch_n8_Vg_global_0_(net1642[0]), .switch_n8_Vg_global_1_(net1641[0]), .switch_n9_Vg_global_0_(net1647[0]), .switch_n9_Vg_global_1_(net1649[0]), .switch_n10_Vg_global_0_(net1647[1]), .switch_n10_Vg_global_1_(net1649[1]), .switch_n11_Vg_global_0_(net1647[2]), .switch_n11_Vg_global_1_(net1649[2]), .switch_n12_Vg_global_0_(net1647[3]), .switch_n12_Vg_global_1_(net1649[3]), .switch_n13_Vg_global_0_(net1647[4]), .switch_n13_Vg_global_1_(net1649[4]), .switch_n14_Vg_global_0_(net1647[5]), .switch_n14_Vg_global_1_(net1649[5]), .switch_n0_VTUN(net1600[0]), .switch_n1_VTUN(net1600[1]), .switch_n2_VTUN(net1600[2]), .switch_n3_VTUN(net1600[3]), .switch_n4_VTUN(net1600[4]), .switch_n5_VTUN(net1600[5]), .switch_n6_VTUN(net1623[0]), .switch_n7_VTUN(net1630[0]), .switch_n8_VTUN(net1637[0]), .switch_n9_VTUN(net1643[0]), .switch_n10_VTUN(net1643[1]), .switch_n11_VTUN(net1643[2]), .switch_n12_VTUN(net1643[3]), .switch_n13_VTUN(net1643[4]), .switch_n14_VTUN(net1643[5]), .switch_n0_VINJ(net1612[0]), .switch_n1_VINJ(net1612[1]), .switch_n2_VINJ(net1612[2]), .switch_n3_VINJ(net1612[3]), .switch_n4_VINJ(net1612[4]), .switch_n5_VINJ(net1612[5]), .switch_n6_VINJ(net1622[0]), .switch_n7_VINJ(net1629[0]), .switch_n8_VINJ(net1636[0]), .switch_n9_VINJ(net1644[0]), .switch_n10_VINJ(net1644[1]), .switch_n11_VINJ(net1644[2]), .switch_n12_VINJ(net1644[3]), .switch_n13_VINJ(net1644[4]), .switch_n14_VINJ(net1644[5]), .switch_n0_Vgrun_r(net1965), .switch_n0_Vgrun(net1877), .switch_n0_AVDD_r(net1969[0]), .switch_n0_run_r(net1872), .switch_n0_prog_r(net1873), .switch_n0_run(net1935));
	none switch_ind(.island_num(1), .direction(horizontal), .col(14));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(15), .VPWR_0_(net1913[0]), .VPWR_1_(net1913[0]), .RUN_IN_0_(net1965), .RUN_IN_1_(net1965), .GND_T(net1645[5]), .VTUN_T(net1643[5]), .decode_0_(net1646[5]), .decode_1_(net1648[5]), .VINJ_T(net1644[5]), .GND(net1535), .CTRL_B_0_(net1533), .prog_r(net1934[0]), .Vg_0_(net1532), .VTUN(net1531), .VINJ(net1534), .VDD_1_(net1969[0]), .PROG(net1873), .RUN(net1872), .Vgsel(net1936));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net903[0:6]), .out_1_row_0(net904[0:6]), .VINJ_0_row_0(net907[0:6]), .VINJ_1_row_0(net908[0:6]), .Vsel_0_row_0(net911[0:6]), .Vsel_1_row_0(net912[0:6]), .Vg_0_row_0(net915[0:6]), .Vg_1_row_0(net916[0:6]), .GNDrow_0(net893[0:6]), .VTUNrow_0(net919[0:6]), .Dcol_0(net112[5:6]), .CLKcol_0(net113[5:6]), .Qcol_5(net236[3:4]), .comcol_0(net1855[0:1]), .VDDcol_0(net1969[0:1]), .Vd_Pcol_0(net1869[0:1]), .Vd_in_0_col_0(net1856[0:1]), .Vd_in_1_col_0(net1860[0:1]), .Vd_in_2_col_0(net1864[0:1]), .Vd_in_3_col_0(net1868[0:1]), .Vd_in_4_col_0(net1857[0:1]), .Vd_in_5_col_0(net1861[0:1]), .Vd_in_6_col_0(net1865[0:1]), .Vd_in_7_col_0(net1869[0:1]), .Vd_o_0_col_5(net1387[0:1]), .Vd_o_1_col_5(net1388[0:1]), .Vd_o_2_col_5(net1389[0:1]), .Vd_o_3_col_5(net1390[0:1]), .Vd_o_4_col_5(net1391[0:1]), .Vd_o_5_col_5(net1392[0:1]), .Vd_o_6_col_5(net1393[0:1]), .Vd_o_7_col_5(net1394[0:1]));

 	/*Programming Mux */ 


	/* Frame */ 
	tile_analog_frame cab_frame(.pin_layer(METAL3), .N_n_gateEN(net1902), .N_n_programdrain(net1903), .N_n_rundrain(net1904), .N_n_cew0(net1878[0]), .N_n_cew1(net1879[0]), .N_n_cew2(net1880[0]), .N_n_cew3(net1881[0]), .N_n_vtun(net1966[0]), .N_n_vinj_0_(net1909), .N_n_vinj_1_(net1910), .N_n_vinj_2_(net1644[5]), .N_n_gnd_0_(net1911), .N_n_gnd_1_(net1912), .N_n_gnd_2_(net1645[5]), .N_n_avdd(net1913[0]), .N_n_s0(net1882[0]), .N_n_s1(net1883[0]), .N_n_s2(net1884[0]), .N_n_s3(net1885[0]), .N_n_s4(net1886[0]), .N_n_s5(net1887[0]), .N_n_s6(net1888[0]), .N_n_s7(net1889[0]), .N_n_s8(net1890[0]), .N_n_s9(net1891[0]), .N_n_s10(net1892[0]), .N_n_s11(net1893[0]), .N_n_s12(net1894), .N_n_s13(net1895), .N_n_s14(net1896), .N_n_s15(net1897), .N_n_s16(net1898), .N_n_s17(net1899), .N_n_s18(net1900), .N_n_s19(net1901), .N_n_prog(net1934[0]), .N_n_run(net1935), .N_n_vgsel(net1936), .S_s_gateEN(net1902), .S_s_programdrain(net1903), .S_s_rundrain(net1904), .S_s_cew0(net1905[0]), .S_s_cew1(net1906[0]), .S_s_cew2(net1907[0]), .S_s_cew3(net1908[0]), .S_s_vtun(net1966[0]), .S_s_vinj_0_(net1909), .S_s_vinj_1_(net1910), .S_s_vinj_2_(net1644[5]), .S_s_gnd_0_(net1911), .S_s_gnd_1_(net1912), .S_s_gnd_2_(net1645[5]), .S_s_avdd(net1913[0]), .S_s_s0(net1914), .S_s_s1(net1915), .S_s_s2(net1916), .S_s_s3(net1917), .S_s_s4(net1918), .S_s_s5(net1919), .S_s_s6(net1920), .S_s_s7(net1921), .S_s_s8(net1922[0]), .S_s_s9(net1923[0]), .S_s_s10(net1924[0]), .S_s_s11(net1925[0]), .S_s_s12(net1926[0]), .S_s_s13(net1927[0]), .S_s_s14(net1928[0]), .S_s_s15(net1929[0]), .S_s_s16(net1930[0]), .S_s_s17(net1931[0]), .S_s_s18(net1932[0]), .S_s_s19(net1933[0]), .S_s_prog(net1934[0]), .S_s_run(net1935), .S_s_vgsel(net1936), .W_w_cns0(net1905[1]), .W_w_cns1(net1906[1]), .W_w_cns2(net1907[1]), .W_w_cns3(net1908[1]), .W_w_vgrun(net1965), .W_w_vtun(net1966[0]), .W_w_vinj(net1644[5]), .W_w_gnd(net1645[5]), .W_w_avdd(net1969[0]), .W_w_drainbit4(net1970), .W_w_drainbit3(net1971), .W_w_drainbit2(net1972), .W_w_drainbit1(net1973), .W_w_drainbit0(net1974), .W_w_s0(net1941[0]), .W_w_s1(net1942[0]), .W_w_s2(net1943[0]), .W_w_s3(net1944[0]), .W_w_s4(net1941[1]), .W_w_s5(net1942[1]), .W_w_s6(net1943[1]), .W_w_s7(net1944[1]), .W_w_s8(net1941[2]), .W_w_s9(net1942[2]), .W_w_s10(net1943[2]), .W_w_s11(net1944[2]), .W_w_s12(net1941[3]), .W_w_s13(net1942[3]), .W_w_s14(net1943[3]), .W_w_s15(net1944[3]), .W_w_s16(net1941[4]), .W_w_s17(net1942[4]), .W_w_s18(net1943[4]), .W_w_s19(net1944[4]), .W_w_drainbit9(net1995), .W_w_drainbit8(net1996), .W_w_drainbit7(net1997), .W_w_drainbit6(net1998), .W_w_drainbit5(net1999), .W_w_drainEN(net2000), .E_e_cns0(net1961[0]), .E_e_cns1(net1962[0]), .E_e_cns2(net1963[0]), .E_e_cns3(net1964[0]), .E_e_vgrun(net1965), .E_e_vtun(net1966[0]), .E_e_vinj(net1644[5]), .E_e_gnd(net1645[5]), .E_e_avdd(net1969[0]), .E_e_drainbit4(net1970), .E_e_drainbit3(net1971), .E_e_drainbit2(net1972), .E_e_drainbit1(net1973), .E_e_drainbit0(net1974), .E_e_s0(net1975[0]), .E_e_s1(net1976[0]), .E_e_s2(net1977[0]), .E_e_s3(net1978[0]), .E_e_s4(net1975[1]), .E_e_s5(net1976[1]), .E_e_s6(net1977[1]), .E_e_s7(net1978[1]), .E_e_s8(net1975[2]), .E_e_s9(net1976[2]), .E_e_s10(net1977[2]), .E_e_s11(net1978[2]), .E_e_s12(net1975[3]), .E_e_s13(net1976[3]), .E_e_s14(net1977[3]), .E_e_s15(net1978[3]), .E_e_s16(net1975[4]), .E_e_s17(net1976[4]), .E_e_s18(net1977[4]), .E_e_s19(net1978[4]), .E_e_drainbit9(net1995), .E_e_drainbit8(net1996), .E_e_drainbit7(net1997), .E_e_drainbit6(net1998), .E_e_drainbit5(net1999), .E_e_drainEN(net2000));
 endmodule