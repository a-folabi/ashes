module TOP(port1);


	/* Island 0 */
	cab1 I__0 (.island_num(0), .row(0), .col(0), .matrix_row(7), .matrix_col(1));
	cab1 I__1 (.island_num(0), .row(0), .col(2), .matrix_row(7), .matrix_col(1));
	cab1 I__2 (.island_num(0), .row(0), .col(4), .matrix_row(7), .matrix_col(1));
	cab1 I__3 (.island_num(0), .row(0), .col(6), .matrix_row(7), .matrix_col(1));
	cab2 I__4 (.island_num(0), .row(0), .col(1), .matrix_row(7), .matrix_col(1));
	cab2 I__5 (.island_num(0), .row(0), .col(3), .matrix_row(7), .matrix_col(1));
	cab2 I__6 (.island_num(0), .row(0), .col(5), .matrix_row(7), .matrix_col(1));

 	/*Programming Mux */ 

 endmodule