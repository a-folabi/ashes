module TOP(port1);


	/* Island 0 */
	TSMC350nm_TA2Cell_Weak I__0 (.island_num(0), .row(0), .col(0), .matrix_row(1), .matrix_col(1), .VIN1_MINUSrow_0(net45), .VIN2_PLUSrow_0(net45), .VIN2_MINUSrow_0(net91), .OUTPUT_0_row_0(net45), .OUTPUT_1_row_0(net45));
	TSMC350nm_TA2Cell_Weak I__1 (.island_num(0), .row(1), .col(0), .matrix_row(1), .matrix_col(1), .VIN1_PLUSrow_0(net45), .VIN1_MINUSrow_0(net91), .VIN2_PLUSrow_0(net91), .VIN2_MINUSrow_0(net46), .OUTPUT_0_row_0(net91), .OUTPUT_1_row_0(net46));
	TSMC350nm_TA2Cell_Weak I__2 (.island_num(0), .row(2), .col(0), .matrix_row(1), .matrix_col(1), .VIN1_PLUSrow_0(net91), .VIN1_MINUSrow_0(net92), .VIN2_PLUSrow_0(net92), .VIN2_MINUSrow_0(net93), .OUTPUT_0_row_0(net92), .OUTPUT_1_row_0(net92));
	TSMC350nm_TA2Cell_Weak I__3 (.island_num(0), .row(3), .col(0), .matrix_row(1), .matrix_col(1), .VIN1_PLUSrow_0(net92), .VIN1_MINUSrow_0(net93), .VIN2_PLUSrow_0(net93), .VIN2_MINUSrow_0(net94), .OUTPUT_0_row_0(net93), .OUTPUT_1_row_0(net94));

 	/*Programming Mux */ 

 endmodule