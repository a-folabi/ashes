module TOP(port1);


	/* Island 0 */
<<<<<<< Updated upstream
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(7), .GND_b_1_row_4(net2030[0:7]), .Vs_b_0_row_4(net124[0:7]), .Vs_b_1_row_4(net125[0:7]), .VINJ_b_1_row_4(net2037[0:7]), .Vsel_b_0_row_4(net1995[0:7]), .Vsel_b_1_row_4(net1996[0:7]), .Vg_b_0_row_4(net2009[0:7]), .Vg_b_1_row_4(net2010[0:7]), .VTUN_brow_4(net2023[0:7]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(17), .matrix_row(5), .matrix_col(9), .GND_b_1_row_4(net2073[0:9]), .Vs_b_0_row_4(net285[0:9]), .Vs_b_1_row_4(net286[0:9]), .VINJ_b_1_row_4(net2072[0:9]), .Vsel_b_0_row_4(net2074[0:9]), .Vsel_b_1_row_4(net2076[0:9]), .Vg_b_0_row_4(net304[0:9]), .Vg_b_1_row_4(net305[0:9]), .VTUN_brow_4(net2071[0:9]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(26), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2050[0:1]), .Vsel_b_0_row_4(net2053[0:1]), .Vsel_b_1_row_4(net2054[0:1]), .Vg_b_0_row_4(net2055[0:1]), .Vg_b_1_row_4(net2056[0:1]), .VTUN_brow_4(net2051[0:1]), .GND_b_1_row_4(net2052[0:1]));
=======
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(0), .matrix_row(5), .matrix_col(7), .GND_b_1_row_4(net2219[0:7]), .Vs_b_0_row_4(net124[0:7]), .Vs_b_1_row_4(net125[0:7]), .VINJ_b_1_row_4(net2226[0:7]), .Vsel_b_0_row_4(net2184[0:7]), .Vsel_b_1_row_4(net2185[0:7]), .Vg_b_0_row_4(net2198[0:7]), .Vg_b_1_row_4(net2199[0:7]), .VTUN_brow_4(net2212[0:7]));
	TSMC350nm_4x2_Indirect I__1 (.island_num(0), .row(0), .col(17), .matrix_row(5), .matrix_col(9), .GND_b_1_row_4(net325[0:9]), .Vs_b_0_row_4(net326[0:9]), .Vs_b_1_row_4(net327[0:9]), .VINJ_b_1_row_4(net345[0:9]), .Vsel_b_0_row_4(net2263[0:9]), .Vsel_b_1_row_4(net2265[0:9]), .Vg_b_0_row_4(net346[0:9]), .Vg_b_1_row_4(net347[0:9]), .VTUN_brow_4(net348[0:9]));
	TSMC350nm_4TGate_ST_BMatrix I__2 (.island_num(0), .row(0), .col(26), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC1_PINS I__3 (.island_num(0), .row(0), .col(7), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2239[0:1]), .Vsel_b_0_row_4(net2242[0:1]), .Vsel_b_1_row_4(net2243[0:1]), .Vg_b_0_row_4(net2244[0:1]), .Vg_b_1_row_4(net2245[0:1]), .VTUN_brow_4(net2240[0:1]), .GND_b_1_row_4(net2241[0:1]));
>>>>>>> Stashed changes
	S_BLOCK_BUFFER I__4 (.island_num(0), .row(0), .col(8), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__5 (.island_num(0), .row(0), .col(9), .matrix_row(4), .matrix_col(1));
	S_BLOCK_CONN_PINS I__6 (.island_num(0), .row(4), .col(9), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__7 (.island_num(0), .row(0), .col(10), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__8 (.island_num(0), .row(3), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__9 (.island_num(0), .row(4), .col(10), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__10 (.island_num(0), .row(0), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_CONN_PINS I__11 (.island_num(0), .row(2), .col(11), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__12 (.island_num(0), .row(3), .col(11), .matrix_row(2), .matrix_col(1));
	S_BLOCK_SPACE_UP_PINS I__13 (.island_num(0), .row(0), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_CONN_PINS I__14 (.island_num(0), .row(1), .col(12), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__15 (.island_num(0), .row(2), .col(12), .matrix_row(3), .matrix_col(1));
	S_BLOCK_CONN_PINS I__16 (.island_num(0), .row(0), .col(13), .matrix_row(1), .matrix_col(1));
	S_BLOCK_SPACE_DOWN_PINS I__17 (.island_num(0), .row(1), .col(13), .matrix_row(4), .matrix_col(1));
<<<<<<< Updated upstream
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2057[0:1]), .Vsel_b_0_row_4(net2060[0:1]), .Vsel_b_1_row_4(net2061[0:1]), .Vg_b_0_row_4(net2062[0:1]), .Vg_b_1_row_4(net2063[0:1]), .VTUN_brow_4(net2058[0:1]), .GND_b_1_row_4(net2059[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2064[0:1]), .Vsel_b_0_row_4(net2067[0:1]), .Vsel_b_1_row_4(net2068[0:1]), .Vg_b_0_row_4(net2069[0:1]), .Vg_b_1_row_4(net2070[0:1]), .VTUN_brow_4(net2065[0:1]), .GND_b_1_row_4(net2066[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(6), .decode_n0_RUN_OUT_0_(net2144), .decode_n0_RUN_OUT_1_(net2145), .decode_n0_RUN_OUT_2_(net2150), .decode_n0_RUN_OUT_3_(net2151), .decode_n1_RUN_OUT_0_(net2156), .decode_n1_RUN_OUT_1_(net2157), .decode_n1_RUN_OUT_2_(net2162), .decode_n1_RUN_OUT_3_(net2163), .decode_n2_RUN_OUT_0_(net2168), .decode_n2_RUN_OUT_1_(net2169), .decode_n2_RUN_OUT_2_(net2174), .decode_n2_RUN_OUT_3_(net2175), .decode_n3_RUN_OUT_0_(net2180), .decode_n3_RUN_OUT_1_(net2181), .decode_n3_RUN_OUT_2_(net2186), .decode_n3_RUN_OUT_3_(net2187), .decode_n4_RUN_OUT_2_(net2192), .decode_n4_RUN_OUT_3_(net2193), .decode_n5_RUN_OUT_0_(net2198), .decode_n5_RUN_OUT_1_(net2199), .decode_n5_RUN_OUT_2_(net2204), .decode_n5_RUN_OUT_3_(net2205), .decode_n6_RUN_OUT_0_(net2210), .decode_n6_RUN_OUT_1_(net2211), .decode_n6_RUN_OUT_2_(net2216), .decode_n6_RUN_OUT_3_(net2217), .decode_n7_RUN_OUT_0_(net2222), .decode_n7_RUN_OUT_1_(net2223), .decode_n7_RUN_OUT_2_(net2228), .decode_n7_RUN_OUT_3_(net2229), .decode_n8_RUN_OUT_0_(net2234), .decode_n8_RUN_OUT_1_(net2235), .decode_n8_RUN_OUT_2_(net2240), .decode_n8_RUN_OUT_3_(net2241), .decode_n9_RUN_OUT_0_(net2246), .decode_n9_RUN_OUT_1_(net2247), .decode_n9_RUN_OUT_2_(net2252), .decode_n9_RUN_OUT_3_(net2253), .decode_n0_OUT_0_(net2142), .decode_n0_OUT_1_(net2143), .decode_n0_OUT_2_(net2148), .decode_n0_OUT_3_(net2149), .decode_n1_OUT_0_(net2154), .decode_n1_OUT_1_(net2155), .decode_n1_OUT_2_(net2160), .decode_n1_OUT_3_(net2161), .decode_n2_OUT_0_(net2166), .decode_n2_OUT_1_(net2167), .decode_n2_OUT_2_(net2172), .decode_n2_OUT_3_(net2173), .decode_n3_OUT_0_(net2178), .decode_n3_OUT_1_(net2179), .decode_n3_OUT_2_(net2184), .decode_n3_OUT_3_(net2185), .decode_n4_OUT_2_(net2190), .decode_n4_OUT_3_(net2191), .decode_n5_OUT_0_(net2196), .decode_n5_OUT_1_(net2197), .decode_n5_OUT_2_(net2202), .decode_n5_OUT_3_(net2203), .decode_n6_OUT_0_(net2208), .decode_n6_OUT_1_(net2209), .decode_n6_OUT_2_(net2214), .decode_n6_OUT_3_(net2215), .decode_n7_OUT_0_(net2220), .decode_n7_OUT_1_(net2221), .decode_n7_OUT_2_(net2226), .decode_n7_OUT_3_(net2227), .decode_n8_OUT_0_(net2232), .decode_n8_OUT_1_(net2233), .decode_n8_OUT_2_(net2238), .decode_n8_OUT_3_(net2239), .decode_n9_OUT_0_(net2244), .decode_n9_OUT_1_(net2245), .decode_n9_OUT_2_(net2250), .decode_n9_OUT_3_(net2251), .decode_n0_VINJ_b_0_(net2140), .decode_n0_VINJ_b_1_(net2146), .decode_n1_VINJ_b_0_(net2152), .decode_n1_VINJ_b_1_(net2158), .decode_n2_VINJ_b_0_(net2164), .decode_n2_VINJ_b_1_(net2170), .decode_n3_VINJ_b_0_(net2176), .decode_n3_VINJ_b_1_(net2182), .decode_n4_VINJ_b_1_(net2188), .decode_n5_VINJ_b_0_(net2194), .decode_n5_VINJ_b_1_(net2200), .decode_n6_VINJ_b_0_(net2206), .decode_n6_VINJ_b_1_(net2212), .decode_n7_VINJ_b_0_(net2218), .decode_n7_VINJ_b_1_(net2224), .decode_n8_VINJ_b_0_(net2230), .decode_n8_VINJ_b_1_(net2236), .decode_n9_VINJ_b_0_(net2242), .decode_n9_VINJ_b_1_(net2248), .decode_n0_GND_b_0_(net2141), .decode_n0_GND_b_1_(net2147), .decode_n1_GND_b_0_(net2153), .decode_n1_GND_b_1_(net2159), .decode_n2_GND_b_0_(net2165), .decode_n2_GND_b_1_(net2171), .decode_n3_GND_b_0_(net2177), .decode_n3_GND_b_1_(net2183), .decode_n4_GND_b_1_(net2189), .decode_n5_GND_b_0_(net2195), .decode_n5_GND_b_1_(net2201), .decode_n6_GND_b_0_(net2207), .decode_n6_GND_b_1_(net2213), .decode_n7_GND_b_0_(net2219), .decode_n7_GND_b_1_(net2225), .decode_n8_GND_b_0_(net2231), .decode_n8_GND_b_1_(net2237), .decode_n9_GND_b_0_(net2243), .decode_n9_GND_b_1_(net2249));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(26), .switch_n0_VPWR_0_(net2144), .switch_n0_VPWR_1_(net2145), .switch_n1_VPWR_0_(net2150), .switch_n1_VPWR_1_(net2151), .switch_n2_VPWR_0_(net2156), .switch_n2_VPWR_1_(net2157), .switch_n3_VPWR_0_(net2162), .switch_n3_VPWR_1_(net2163), .switch_n4_VPWR_0_(net2168), .switch_n4_VPWR_1_(net2169), .switch_n5_VPWR_0_(net2174), .switch_n5_VPWR_1_(net2175), .switch_n6_VPWR_0_(net2180), .switch_n6_VPWR_1_(net2181), .switch_n7_VPWR_0_(net2186), .switch_n7_VPWR_1_(net2187), .switch_n14_VPWR_0_(net2192), .switch_n14_VPWR_1_(net2193), .switch_n16_VPWR_0_(net2198), .switch_n16_VPWR_1_(net2199), .switch_n17_VPWR_0_(net2204), .switch_n17_VPWR_1_(net2205), .switch_n18_VPWR_0_(net2210), .switch_n18_VPWR_1_(net2211), .switch_n19_VPWR_0_(net2216), .switch_n19_VPWR_1_(net2217), .switch_n20_VPWR_0_(net2222), .switch_n20_VPWR_1_(net2223), .switch_n21_VPWR_0_(net2228), .switch_n21_VPWR_1_(net2229), .switch_n22_VPWR_0_(net2234), .switch_n22_VPWR_1_(net2235), .switch_n23_VPWR_0_(net2240), .switch_n23_VPWR_1_(net2241), .switch_n24_VPWR_0_(net2246), .switch_n24_VPWR_1_(net2247), .switch_n25_VPWR_0_(net2252), .switch_n25_VPWR_1_(net2253), .switch_n0_GND_T(net2141), .switch_n1_GND_T(net2147), .switch_n2_GND_T(net2153), .switch_n3_GND_T(net2159), .switch_n4_GND_T(net2165), .switch_n5_GND_T(net2171), .switch_n6_GND_T(net2177), .switch_n7_GND_T(net2183), .switch_n14_GND_T(net2189), .switch_n16_GND_T(net2195), .switch_n17_GND_T(net2201), .switch_n18_GND_T(net2207), .switch_n19_GND_T(net2213), .switch_n20_GND_T(net2219), .switch_n21_GND_T(net2225), .switch_n22_GND_T(net2231), .switch_n23_GND_T(net2237), .switch_n24_GND_T(net2243), .switch_n25_GND_T(net2249), .switch_n0_decode_0_(net2142), .switch_n0_decode_1_(net2143), .switch_n1_decode_0_(net2148), .switch_n1_decode_1_(net2149), .switch_n2_decode_0_(net2154), .switch_n2_decode_1_(net2155), .switch_n3_decode_0_(net2160), .switch_n3_decode_1_(net2161), .switch_n4_decode_0_(net2166), .switch_n4_decode_1_(net2167), .switch_n5_decode_0_(net2172), .switch_n5_decode_1_(net2173), .switch_n6_decode_0_(net2178), .switch_n6_decode_1_(net2179), .switch_n7_decode_0_(net2184), .switch_n7_decode_1_(net2185), .switch_n14_decode_0_(net2190), .switch_n14_decode_1_(net2191), .switch_n16_decode_0_(net2196), .switch_n16_decode_1_(net2197), .switch_n17_decode_0_(net2202), .switch_n17_decode_1_(net2203), .switch_n18_decode_0_(net2208), .switch_n18_decode_1_(net2209), .switch_n19_decode_0_(net2214), .switch_n19_decode_1_(net2215), .switch_n20_decode_0_(net2220), .switch_n20_decode_1_(net2221), .switch_n21_decode_0_(net2226), .switch_n21_decode_1_(net2227), .switch_n22_decode_0_(net2232), .switch_n22_decode_1_(net2233), .switch_n23_decode_0_(net2238), .switch_n23_decode_1_(net2239), .switch_n24_decode_0_(net2244), .switch_n24_decode_1_(net2245), .switch_n25_decode_0_(net2250), .switch_n25_decode_1_(net2251), .switch_n0_VINJ_T(net2140), .switch_n1_VINJ_T(net2146), .switch_n2_VINJ_T(net2152), .switch_n3_VINJ_T(net2158), .switch_n4_VINJ_T(net2164), .switch_n5_VINJ_T(net2170), .switch_n6_VINJ_T(net2176), .switch_n7_VINJ_T(net2182), .switch_n14_VINJ_T(net2188), .switch_n16_VINJ_T(net2194), .switch_n17_VINJ_T(net2200), .switch_n18_VINJ_T(net2206), .switch_n19_VINJ_T(net2212), .switch_n20_VINJ_T(net2218), .switch_n21_VINJ_T(net2224), .switch_n22_VINJ_T(net2230), .switch_n23_VINJ_T(net2236), .switch_n24_VINJ_T(net2242), .switch_n25_VINJ_T(net2248));
=======
	S_BLOCK_SEC2_PINS I__18 (.island_num(0), .row(0), .col(14), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2246[0:1]), .Vsel_b_0_row_4(net2249[0:1]), .Vsel_b_1_row_4(net2250[0:1]), .Vg_b_0_row_4(net2251[0:1]), .Vg_b_1_row_4(net2252[0:1]), .VTUN_brow_4(net2247[0:1]), .GND_b_1_row_4(net2248[0:1]));
	S_BLOCK_23CONN I__19 (.island_num(0), .row(0), .col(15), .matrix_row(5), .matrix_col(1));
	S_BLOCK_SEC3_PINS I__20 (.island_num(0), .row(0), .col(16), .matrix_row(5), .matrix_col(1), .VINJ_brow_4(net2253[0:1]), .Vsel_b_0_row_4(net2256[0:1]), .Vsel_b_1_row_4(net2257[0:1]), .Vg_b_0_row_4(net2258[0:1]), .Vg_b_1_row_4(net2259[0:1]), .VTUN_brow_4(net2254[0:1]), .GND_b_1_row_4(net2255[0:1]));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(6), .decode_n0_RUN_OUT_0_(net2330), .decode_n0_RUN_OUT_1_(net2331), .decode_n0_RUN_OUT_2_(net2336), .decode_n0_RUN_OUT_3_(net2337), .decode_n1_RUN_OUT_0_(net2342), .decode_n1_RUN_OUT_1_(net2343), .decode_n1_RUN_OUT_2_(net2348), .decode_n1_RUN_OUT_3_(net2349), .decode_n2_RUN_OUT_0_(net2354), .decode_n2_RUN_OUT_1_(net2355), .decode_n2_RUN_OUT_2_(net2360), .decode_n2_RUN_OUT_3_(net2361), .decode_n3_RUN_OUT_0_(net2366), .decode_n3_RUN_OUT_1_(net2367), .decode_n3_RUN_OUT_2_(net2372), .decode_n3_RUN_OUT_3_(net2373), .decode_n4_RUN_OUT_2_(net2378), .decode_n4_RUN_OUT_3_(net2379), .decode_n5_RUN_OUT_0_(net2384), .decode_n5_RUN_OUT_1_(net2385), .decode_n5_RUN_OUT_2_(net2390), .decode_n5_RUN_OUT_3_(net2391), .decode_n6_RUN_OUT_0_(net2396), .decode_n6_RUN_OUT_1_(net2397), .decode_n6_RUN_OUT_2_(net2402), .decode_n6_RUN_OUT_3_(net2403), .decode_n7_RUN_OUT_0_(net2408), .decode_n7_RUN_OUT_1_(net2409), .decode_n7_RUN_OUT_2_(net2414), .decode_n7_RUN_OUT_3_(net2415), .decode_n8_RUN_OUT_0_(net2420), .decode_n8_RUN_OUT_1_(net2421), .decode_n8_RUN_OUT_2_(net2426), .decode_n8_RUN_OUT_3_(net2427), .decode_n9_RUN_OUT_0_(net2432), .decode_n9_RUN_OUT_1_(net2433), .decode_n9_RUN_OUT_2_(net2438), .decode_n9_RUN_OUT_3_(net2439), .decode_n0_OUT_0_(net2328), .decode_n0_OUT_1_(net2329), .decode_n0_OUT_2_(net2334), .decode_n0_OUT_3_(net2335), .decode_n1_OUT_0_(net2340), .decode_n1_OUT_1_(net2341), .decode_n1_OUT_2_(net2346), .decode_n1_OUT_3_(net2347), .decode_n2_OUT_0_(net2352), .decode_n2_OUT_1_(net2353), .decode_n2_OUT_2_(net2358), .decode_n2_OUT_3_(net2359), .decode_n3_OUT_0_(net2364), .decode_n3_OUT_1_(net2365), .decode_n3_OUT_2_(net2370), .decode_n3_OUT_3_(net2371), .decode_n4_OUT_2_(net2376), .decode_n4_OUT_3_(net2377), .decode_n5_OUT_0_(net2382), .decode_n5_OUT_1_(net2383), .decode_n5_OUT_2_(net2388), .decode_n5_OUT_3_(net2389), .decode_n6_OUT_0_(net2394), .decode_n6_OUT_1_(net2395), .decode_n6_OUT_2_(net2400), .decode_n6_OUT_3_(net2401), .decode_n7_OUT_0_(net2406), .decode_n7_OUT_1_(net2407), .decode_n7_OUT_2_(net2412), .decode_n7_OUT_3_(net2413), .decode_n8_OUT_0_(net2418), .decode_n8_OUT_1_(net2419), .decode_n8_OUT_2_(net2424), .decode_n8_OUT_3_(net2425), .decode_n9_OUT_0_(net2430), .decode_n9_OUT_1_(net2431), .decode_n9_OUT_2_(net2436), .decode_n9_OUT_3_(net2437), .decode_n0_VINJ_b_0_(net2326), .decode_n0_VINJ_b_1_(net2332), .decode_n1_VINJ_b_0_(net2338), .decode_n1_VINJ_b_1_(net2344), .decode_n2_VINJ_b_0_(net2350), .decode_n2_VINJ_b_1_(net2356), .decode_n3_VINJ_b_0_(net2362), .decode_n3_VINJ_b_1_(net2368), .decode_n4_VINJ_b_1_(net2374), .decode_n5_VINJ_b_0_(net2380), .decode_n5_VINJ_b_1_(net2386), .decode_n6_VINJ_b_0_(net2392), .decode_n6_VINJ_b_1_(net2398), .decode_n7_VINJ_b_0_(net2404), .decode_n7_VINJ_b_1_(net2410), .decode_n8_VINJ_b_0_(net2416), .decode_n8_VINJ_b_1_(net2422), .decode_n9_VINJ_b_0_(net2428), .decode_n9_VINJ_b_1_(net2434), .decode_n0_GND_b_0_(net2327), .decode_n0_GND_b_1_(net2333), .decode_n1_GND_b_0_(net2339), .decode_n1_GND_b_1_(net2345), .decode_n2_GND_b_0_(net2351), .decode_n2_GND_b_1_(net2357), .decode_n3_GND_b_0_(net2363), .decode_n3_GND_b_1_(net2369), .decode_n4_GND_b_1_(net2375), .decode_n5_GND_b_0_(net2381), .decode_n5_GND_b_1_(net2387), .decode_n6_GND_b_0_(net2393), .decode_n6_GND_b_1_(net2399), .decode_n7_GND_b_0_(net2405), .decode_n7_GND_b_1_(net2411), .decode_n8_GND_b_0_(net2417), .decode_n8_GND_b_1_(net2423), .decode_n9_GND_b_0_(net2429), .decode_n9_GND_b_1_(net2435));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(26), .switch_n0_VPWR_0_(net2330), .switch_n0_VPWR_1_(net2331), .switch_n1_VPWR_0_(net2336), .switch_n1_VPWR_1_(net2337), .switch_n2_VPWR_0_(net2342), .switch_n2_VPWR_1_(net2343), .switch_n3_VPWR_0_(net2348), .switch_n3_VPWR_1_(net2349), .switch_n4_VPWR_0_(net2354), .switch_n4_VPWR_1_(net2355), .switch_n5_VPWR_0_(net2360), .switch_n5_VPWR_1_(net2361), .switch_n6_VPWR_0_(net2366), .switch_n6_VPWR_1_(net2367), .switch_n7_VPWR_0_(net2372), .switch_n7_VPWR_1_(net2373), .switch_n14_VPWR_0_(net2378), .switch_n14_VPWR_1_(net2379), .switch_n16_VPWR_0_(net2384), .switch_n16_VPWR_1_(net2385), .switch_n17_VPWR_0_(net2390), .switch_n17_VPWR_1_(net2391), .switch_n18_VPWR_0_(net2396), .switch_n18_VPWR_1_(net2397), .switch_n19_VPWR_0_(net2402), .switch_n19_VPWR_1_(net2403), .switch_n20_VPWR_0_(net2408), .switch_n20_VPWR_1_(net2409), .switch_n21_VPWR_0_(net2414), .switch_n21_VPWR_1_(net2415), .switch_n22_VPWR_0_(net2420), .switch_n22_VPWR_1_(net2421), .switch_n23_VPWR_0_(net2426), .switch_n23_VPWR_1_(net2427), .switch_n24_VPWR_0_(net2432), .switch_n24_VPWR_1_(net2433), .switch_n25_VPWR_0_(net2438), .switch_n25_VPWR_1_(net2439), .switch_n0_GND_T(net2327), .switch_n1_GND_T(net2333), .switch_n2_GND_T(net2339), .switch_n3_GND_T(net2345), .switch_n4_GND_T(net2351), .switch_n5_GND_T(net2357), .switch_n6_GND_T(net2363), .switch_n7_GND_T(net2369), .switch_n14_GND_T(net2375), .switch_n16_GND_T(net2381), .switch_n17_GND_T(net2387), .switch_n18_GND_T(net2393), .switch_n19_GND_T(net2399), .switch_n20_GND_T(net2405), .switch_n21_GND_T(net2411), .switch_n22_GND_T(net2417), .switch_n23_GND_T(net2423), .switch_n24_GND_T(net2429), .switch_n25_GND_T(net2435), .switch_n0_decode_0_(net2328), .switch_n0_decode_1_(net2329), .switch_n1_decode_0_(net2334), .switch_n1_decode_1_(net2335), .switch_n2_decode_0_(net2340), .switch_n2_decode_1_(net2341), .switch_n3_decode_0_(net2346), .switch_n3_decode_1_(net2347), .switch_n4_decode_0_(net2352), .switch_n4_decode_1_(net2353), .switch_n5_decode_0_(net2358), .switch_n5_decode_1_(net2359), .switch_n6_decode_0_(net2364), .switch_n6_decode_1_(net2365), .switch_n7_decode_0_(net2370), .switch_n7_decode_1_(net2371), .switch_n14_decode_0_(net2376), .switch_n14_decode_1_(net2377), .switch_n16_decode_0_(net2382), .switch_n16_decode_1_(net2383), .switch_n17_decode_0_(net2388), .switch_n17_decode_1_(net2389), .switch_n18_decode_0_(net2394), .switch_n18_decode_1_(net2395), .switch_n19_decode_0_(net2400), .switch_n19_decode_1_(net2401), .switch_n20_decode_0_(net2406), .switch_n20_decode_1_(net2407), .switch_n21_decode_0_(net2412), .switch_n21_decode_1_(net2413), .switch_n22_decode_0_(net2418), .switch_n22_decode_1_(net2419), .switch_n23_decode_0_(net2424), .switch_n23_decode_1_(net2425), .switch_n24_decode_0_(net2430), .switch_n24_decode_1_(net2431), .switch_n25_decode_0_(net2436), .switch_n25_decode_1_(net2437), .switch_n0_VINJ_T(net2326), .switch_n1_VINJ_T(net2332), .switch_n2_VINJ_T(net2338), .switch_n3_VINJ_T(net2344), .switch_n4_VINJ_T(net2350), .switch_n5_VINJ_T(net2356), .switch_n6_VINJ_T(net2362), .switch_n7_VINJ_T(net2368), .switch_n14_VINJ_T(net2374), .switch_n16_VINJ_T(net2380), .switch_n17_VINJ_T(net2386), .switch_n18_VINJ_T(net2392), .switch_n19_VINJ_T(net2398), .switch_n20_VINJ_T(net2404), .switch_n21_VINJ_T(net2410), .switch_n22_VINJ_T(net2416), .switch_n23_VINJ_T(net2422), .switch_n24_VINJ_T(net2428), .switch_n25_VINJ_T(net2434));
>>>>>>> Stashed changes
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch));
	none switch_ind(.island_num(0), .direction(horizontal), .col(8));
	none switch_ind(.island_num(0), .direction(horizontal), .col(9));
	none switch_ind(.island_num(0), .direction(horizontal), .col(10));
	none switch_ind(.island_num(0), .direction(horizontal), .col(11));
	none switch_ind(.island_num(0), .direction(horizontal), .col(12));
	none switch_ind(.island_num(0), .direction(horizontal), .col(13));
	none switch_ind(.island_num(0), .direction(horizontal), .col(15));


	/* Island 1 */
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__0 (.island_num(1), .row(0), .col(0), .matrix_row(1), .matrix_col(8));
<<<<<<< Updated upstream
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(7), .matrix_col(8), .GND_b_0_row_6(net1138[0:8]), .GND_b_1_row_6(net1139[0:8]), .Vs_b_0_row_6(net1148[0:8]), .Vs_b_1_row_6(net1149[0:8]), .VINJ_b_0_row_6(net1152[0:8]), .VINJ_b_1_row_6(net1153[0:8]), .Vsel_b_0_row_6(net1156[0:8]), .Vsel_b_1_row_6(net1157[0:8]), .Vg_b_0_row_6(net1160[0:8]), .Vg_b_1_row_6(net1161[0:8]), .VTUN_brow_6(net1164[0:8]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(8), .matrix_row(6), .matrix_col(10));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(7), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1895), .P_1_row_0(net1896), .A_0_row_0(net1897), .A_1_row_0(net1898), .A_2_row_0(net1899), .A_3_row_0(net1900));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1908), .P_1_row_0(net1909), .A_0_row_0(net1910), .A_1_row_0(net1911), .A_2_row_0(net1912), .A_3_row_0(net1913));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1926), .P_1_row_0(net1927), .A_0_row_0(net1928), .A_1_row_0(net1929), .A_2_row_0(net1930), .A_3_row_0(net1931));
	TSMC350nm_4TGate_ST_BMatrix_NoSwitch I__8 (.island_num(1), .row(3), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1944), .P_1_row_0(net1945), .P_2_row_0(net1946), .P_3_row_0(net1947), .A_0_row_0(net1948), .A_1_row_0(net1949), .A_2_row_0(net1950), .A_3_row_0(net1951));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net1963), .P_1_row_0(net1964), .P_2_row_0(net1965), .P_3_row_0(net1966), .A_0_row_0(net1967), .A_1_row_0(net1968));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1978), .A_1_row_0(net1979), .A_2_row_0(net1980), .A_3_row_0(net1981));
	TSMC350nm_4TGate_ST_BMatrix I__11 (.island_num(1), .row(6), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net1985), .A_1_row_0(net1986), .A_2_row_0(net1987), .A_3_row_0(net1988));
=======
	TSMC350nm_4x2_Indirect I__1 (.island_num(1), .row(1), .col(0), .matrix_row(7), .matrix_col(8), .GND_b_0_row_6(net1221[0:8]), .GND_b_1_row_6(net1222[0:8]), .Vs_b_0_row_6(net1231[0:8]), .Vs_b_1_row_6(net1232[0:8]), .VINJ_b_0_row_6(net1235[0:8]), .VINJ_b_1_row_6(net1236[0:8]), .Vsel_b_0_row_6(net1239[0:8]), .Vsel_b_1_row_6(net1240[0:8]), .Vg_b_0_row_6(net1243[0:8]), .Vg_b_1_row_6(net1244[0:8]), .VTUN_brow_6(net1247[0:8]));
	TSMC350nm_4x2_Indirect_top_AorB_matrx I__2 (.island_num(1), .row(0), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__3 (.island_num(1), .row(1), .col(8), .matrix_row(6), .matrix_col(10));
	TSMC350nm_4x2_Indirect_bot_B_matrx I__4 (.island_num(1), .row(7), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4TGate_ST_BMatrix I__5 (.island_num(1), .row(0), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2083), .P_1_row_0(net2084), .A_0_row_0(net2085), .A_1_row_0(net2086), .A_2_row_0(net2087), .A_3_row_0(net2088));
	TSMC350nm_4TGate_ST_BMatrix I__6 (.island_num(1), .row(1), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2096), .P_1_row_0(net2097), .A_0_row_0(net2098), .A_1_row_0(net2099), .A_2_row_0(net2100), .A_3_row_0(net2101));
	TSMC350nm_4TGate_ST_BMatrix I__7 (.island_num(1), .row(2), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2114), .P_1_row_0(net2115), .A_0_row_0(net2116), .A_1_row_0(net2117), .A_2_row_0(net2118), .A_3_row_0(net2119));
	TSMC350nm_4TGate_ST_BMatrix_NoSwitch I__8 (.island_num(1), .row(3), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2132), .P_1_row_0(net2133), .P_2_row_0(net2134), .P_3_row_0(net2135), .A_0_row_0(net2136), .A_1_row_0(net2137), .A_2_row_0(net2138), .A_3_row_0(net2139));
	TSMC350nm_4TGate_ST_BMatrix I__9 (.island_num(1), .row(4), .col(18), .matrix_row(1), .matrix_col(1), .P_0_row_0(net2151), .P_1_row_0(net2152), .P_2_row_0(net2153), .P_3_row_0(net2154), .A_0_row_0(net2155), .A_1_row_0(net2156));
	TSMC350nm_4TGate_ST_BMatrix I__10 (.island_num(1), .row(5), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net2166), .A_1_row_0(net2167), .A_2_row_0(net2168), .A_3_row_0(net2169));
	TSMC350nm_4TGate_ST_BMatrix I__11 (.island_num(1), .row(6), .col(18), .matrix_row(1), .matrix_col(1), .A_0_row_0(net2174), .A_1_row_0(net2175), .A_2_row_0(net2176), .A_3_row_0(net2177));
>>>>>>> Stashed changes
	TSMC350nm_4TGate_ST_BMatrix I__12 (.island_num(1), .row(7), .col(18), .matrix_row(1), .matrix_col(1));
	TSMC350nm_OutMtrx_IndrctSwcs I__13 (.island_num(1), .row(9), .col(8), .matrix_row(1), .matrix_col(10));
	TSMC350nm_4x2_Indirect I__14 (.island_num(1), .row(10), .col(8), .matrix_row(2), .matrix_col(10), .Vd_Rl_0_col_0(net1917[0:2]), .Vd_Rl_1_col_0(net1918[0:2]), .Vd_Rl_2_col_0(net1919[0:2]), .Vd_Rl_3_col_0(net1920[0:2]), .Vd_Pl_0_col_0(net1921[0:2]), .Vd_Pl_1_col_0(net1922[0:2]), .Vd_Pl_2_col_0(net1923[0:2]), .Vd_Pl_3_col_0(net1924[0:2]));
	TSMC350nm_4TGate_ST_BMatrix I__15 (.island_num(1), .row(10), .col(18), .matrix_row(2), .matrix_col(1));
<<<<<<< Updated upstream
	TSMC350nm_TA2Cell_Weak cab_device_16 (.island_num(1), .row(2), .col(19), .VD_P_0_(net1895), .VD_P_1_(net1896), .VIN1_PLUS(net1897), .VIN1_MINUS(net1898), .VIN2_PLUS(net1899), .VIN2_MINUS(net1900), .OUTPUT_0_(net1901[0]), .OUTPUT_1_(net1902[0]), .Vsel_0_(net1972), .Vsel_1_(net1973), .RUN(net1903), .Vg_0_(net1974), .Vg_1_(net1975), .PROG(net1904), .VTUN(net1905), .VINJ(net1906), .GND(net1907), .VPWR(net2317[0]), .Vsel_b_0_(net1916), .Vsel_b_1_(net1917), .RUN_b(net1918), .Vg_b_0_(net1919), .Vg_b_1_(net1920), .PROG_b(net1921), .VTUN_b(net1922), .VINJ_b(net1923), .GND_b(net1924), .VPWR_b(net1925));
	TSMC350nm_TA2Cell_Weak cab_device_17 (.island_num(1), .row(3), .col(19), .VD_P_0_(net1908), .VD_P_1_(net1909), .VIN1_PLUS(net1910), .VIN1_MINUS(net1911), .VIN2_PLUS(net1912), .VIN2_MINUS(net1913), .OUTPUT_0_(net1914[0]), .OUTPUT_1_(net1915[0]), .Vsel_0_(net1916), .Vsel_1_(net1917), .RUN(net1918), .Vg_0_(net1919), .Vg_1_(net1920), .PROG(net1921), .VTUN(net1922), .VINJ(net1923), .GND(net1924), .VPWR(net1925), .Vsel_b_0_(net1934), .Vsel_b_1_(net1935), .RUN_b(net1936), .Vg_b_0_(net1937), .Vg_b_1_(net1938), .PROG_b(net1939), .VTUN_b(net1940), .VINJ_b(net1941), .GND_b(net1942), .VPWR_b(net1943));
	TSMC350nm_TA2Cell_Strong cab_device_18 (.island_num(1), .row(4), .col(19), .VD_P_0_(net1926), .VD_P_1_(net1927), .VIN1_PLUS(net1928), .VIN1_MINUS(net1929), .VIN2_PLUS(net1930), .VIN2_MINUS(net1931), .OUTPUT_0_(net1932[0]), .OUTPUT_1_(net1933[0]), .Vsel_0_(net1934), .Vsel_1_(net1935), .RUN(net1936), .Vg_0_(net1937), .Vg_1_(net1938), .PROG(net1939), .VTUN(net1940), .VINJ(net1941), .GND(net1942), .VPWR(net1943), .Vg_b_0_(net1959), .PROG_b(net1962), .VTUN_b(net1960), .VINJ_b(net1958), .GND_b(net1961));
	TSMC350nm_4WTA_IndirectProg cab_device_19 (.island_num(1), .row(5), .col(19), .VD_P_0_(net1944), .VD_P_1_(net1945), .VD_P_2_(net1946), .VD_P_3_(net1947), .Iin_0_(net1948), .Iin_1_(net1949), .Iin_2_(net1950), .Iin_3_(net1951), .Vout_0_(net1952[0]), .Vout_1_(net1953[0]), .Vout_2_(net1954[0]), .Vout_3_(net1955[0]), .Vmid(net1956[0]), .Vbias(net1957[0]), .Vsel(net1972), .Vs(net2317[0]), .VINJ(net1958), .Vg(net1959), .VTUN(net1960), .GND(net1961), .PROG(net1962), .VINJ_b(net1971), .VTUN_b(net1977), .GND_b(net1976));
	TSMC350nm_Cap_Bank cab_device_20 (.island_num(1), .row(6), .col(19), .VD_P_0_(net1963), .VD_P_1_(net1964), .VD_P_2_(net1965), .VD_P_3_(net1966), .VIN_0_(net1967), .VIN_1_(net1968), .OUT_0_(net1969[0]), .OUT_1_(net1970[0]), .VINJ(net1971), .Vsel_0_(net1972), .Vsel_1_(net1973), .Vg_0_(net1974), .Vg_1_(net1975), .GND(net1976), .VTUN(net1977), .GND_b(net1984));
	TSMC350nm_NandPfets cab_device_21 (.island_num(1), .row(7), .col(19), .GATE_N(net1978), .SOURCE_N(net1979), .GATE_P(net1980), .SOURCE_P(net1981), .DRAIN_N(net1982[0]), .DRAIN_P(net1983[0]), .VPWR(net2317[0]), .GND(net1984), .VPWR_b(net1992), .GND_b(net1993));
	TSMC350nm_TGate_2nMirror cab_device_22 (.island_num(1), .row(8), .col(19), .IN_CM_0_(net1985), .IN_CM_1_(net1986), .SelN(net1987), .IN_TG(net1988), .OUT_CM_0_(net1989[0]), .OUT_CM_1_(net1990[0]), .OUT_TG(net1991[0]), .VPWR(net1992), .GND(net1993));
=======
	TSMC350nm_TA2Cell_Weak cab_device_16 (.island_num(1), .row(2), .col(19), .VD_P_0_(net2083), .VD_P_1_(net2084), .VIN1_PLUS(net2085), .VIN1_MINUS(net2086), .VIN2_PLUS(net2087), .VIN2_MINUS(net2088), .OUTPUT_0_(net2089[0]), .OUTPUT_1_(net2090[0]), .Vsel_0_(net2160), .Vsel_1_(net2161), .RUN(net2091), .Vg_0_(net2162), .Vg_1_(net2163), .PROG(net2092), .VTUN(net2093), .VINJ(net2094), .GND(net2095), .VPWR(net2172), .Vsel_b_0_(net2104), .Vsel_b_1_(net2105), .RUN_b(net2106), .Vg_b_0_(net2107), .Vg_b_1_(net2108), .PROG_b(net2109), .VTUN_b(net2110), .VINJ_b(net2111), .GND_b(net2112), .VPWR_b(net2113));
	TSMC350nm_TA2Cell_Weak cab_device_17 (.island_num(1), .row(3), .col(19), .VD_P_0_(net2096), .VD_P_1_(net2097), .VIN1_PLUS(net2098), .VIN1_MINUS(net2099), .VIN2_PLUS(net2100), .VIN2_MINUS(net2101), .OUTPUT_0_(net2102[0]), .OUTPUT_1_(net2103[0]), .Vsel_0_(net2104), .Vsel_1_(net2105), .RUN(net2106), .Vg_0_(net2107), .Vg_1_(net2108), .PROG(net2109), .VTUN(net2110), .VINJ(net2111), .GND(net2112), .VPWR(net2113), .Vsel_b_0_(net2122), .Vsel_b_1_(net2123), .RUN_b(net2124), .Vg_b_0_(net2125), .Vg_b_1_(net2126), .PROG_b(net2127), .VTUN_b(net2128), .VINJ_b(net2129), .GND_b(net2130), .VPWR_b(net2131));
	TSMC350nm_TA2Cell_Strong cab_device_18 (.island_num(1), .row(4), .col(19), .VD_P_0_(net2114), .VD_P_1_(net2115), .VIN1_PLUS(net2116), .VIN1_MINUS(net2117), .VIN2_PLUS(net2118), .VIN2_MINUS(net2119), .OUTPUT_0_(net2120[0]), .OUTPUT_1_(net2121[0]), .Vsel_0_(net2122), .Vsel_1_(net2123), .RUN(net2124), .Vg_0_(net2125), .Vg_1_(net2126), .PROG(net2127), .VTUN(net2128), .VINJ(net2129), .GND(net2130), .VPWR(net2131), .Vg_b_0_(net2147), .PROG_b(net2150), .VTUN_b(net2148), .VINJ_b(net2146), .GND_b(net2149));
	TSMC350nm_4WTA_IndirectProg cab_device_19 (.island_num(1), .row(5), .col(19), .VD_P_0_(net2132), .VD_P_1_(net2133), .VD_P_2_(net2134), .VD_P_3_(net2135), .Iin_0_(net2136), .Iin_1_(net2137), .Iin_2_(net2138), .Iin_3_(net2139), .Vout_0_(net2140[0]), .Vout_1_(net2141[0]), .Vout_2_(net2142[0]), .Vout_3_(net2143[0]), .Vmid(net2144[0]), .Vbias(net2145[0]), .Vsel(net2160), .Vs(net2172), .VINJ(net2146), .Vg(net2147), .VTUN(net2148), .GND(net2149), .PROG(net2150), .VINJ_b(net2159), .VTUN_b(net2165), .GND_b(net2164));
	TSMC350nm_Cap_Bank cab_device_20 (.island_num(1), .row(6), .col(19), .VD_P_0_(net2151), .VD_P_1_(net2152), .VD_P_2_(net2153), .VD_P_3_(net2154), .VIN_0_(net2155), .VIN_1_(net2156), .OUT_0_(net2157[0]), .OUT_1_(net2158[0]), .VINJ(net2159), .Vsel_0_(net2160), .Vsel_1_(net2161), .Vg_0_(net2162), .Vg_1_(net2163), .GND(net2164), .VTUN(net2165), .GND_b(net2173));
	TSMC350nm_NandPfets cab_device_21 (.island_num(1), .row(7), .col(19), .GATE_N(net2166), .SOURCE_N(net2167), .GATE_P(net2168), .SOURCE_P(net2169), .DRAIN_N(net2170[0]), .DRAIN_P(net2171[0]), .VPWR(net2172), .GND(net2173), .VPWR_b(net2181), .GND_b(net2182));
	TSMC350nm_TGate_2nMirror cab_device_22 (.island_num(1), .row(8), .col(19), .IN_CM_0_(net2174), .IN_CM_1_(net2175), .SelN(net2176), .IN_TG(net2177), .OUT_CM_0_(net2178[0]), .OUT_CM_1_(net2179[0]), .OUT_TG(net2180[0]), .VPWR(net2181), .GND(net2182));
>>>>>>> Stashed changes

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(1), .direction(vertical), .bits(6));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(1), .direction(vertical), .num(12), .type(drain_select));
<<<<<<< Updated upstream
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(12), .type(prog_switch), .switch_n8_PR_3_(net2318[0]));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(20), .switch_n0_Input_0_(net1994), .switch_n0_Input_1_(net2030[0]), .switch_n1_Input_0_(net124[1]), .switch_n1_Input_1_(net125[1]), .switch_n2_Input_0_(net124[2]), .switch_n2_Input_1_(net125[2]), .switch_n3_Input_0_(net124[3]), .switch_n3_Input_1_(net125[3]), .switch_n4_Input_0_(net285[0]), .switch_n4_Input_1_(net286[0]), .switch_n5_Input_0_(net285[1]), .switch_n5_Input_1_(net286[1]), .switch_n6_Input_0_(net285[2]), .switch_n6_Input_1_(net286[2]), .switch_n7_Input_0_(net285[3]), .switch_n7_Input_1_(net286[3]), .switch_n8_Input_0_(net2316[0]), .switch_n8_Input_1_(net1901[0]), .switch_n9_Input_0_(net1902[0]), .switch_n9_Input_1_(net1914[0]), .switch_n10_Input_0_(net1915[0]), .switch_n10_Input_1_(net1932[0]), .switch_n11_Input_0_(net1933[0]), .switch_n11_Input_1_(net1952[0]), .switch_n12_Input_0_(net1953[0]), .switch_n12_Input_1_(net1954[0]), .switch_n13_Input_0_(net1955[0]), .switch_n13_Input_1_(net1956[0]), .switch_n14_Input_0_(net1957[0]), .switch_n14_Input_1_(net1969[0]), .switch_n15_Input_0_(net1970[0]), .switch_n15_Input_1_(net1982[0]), .switch_n16_Input_0_(net1983[0]), .switch_n16_Input_1_(net1989[0]), .switch_n17_Input_0_(net1990[0]), .switch_n17_Input_1_(net1991[0]), .switch_n0_GND(net2030[0]), .switch_n1_GND(net2030[1]), .switch_n2_GND(net2030[2]), .switch_n3_GND(net2030[3]), .switch_n4_GND(net2030[4]), .switch_n5_GND(net2030[5]), .switch_n6_GND(net2030[6]), .switch_n7_GND(net2052[0]), .switch_n8_GND(net2059[0]), .switch_n9_GND(net2066[0]), .switch_n10_GND(net2073[0]), .switch_n11_GND(net2073[1]), .switch_n12_GND(net2073[2]), .switch_n13_GND(net2073[3]), .switch_n14_GND(net2073[4]), .switch_n15_GND(net2073[5]), .switch_n16_GND(net2073[6]), .switch_n17_GND(net2073[7]), .switch_n0_Vsel_0_(net1995[0]), .switch_n0_Vsel_1_(net1996[0]), .switch_n1_Vsel_0_(net1995[1]), .switch_n1_Vsel_1_(net1996[1]), .switch_n2_Vsel_0_(net1995[2]), .switch_n2_Vsel_1_(net1996[2]), .switch_n3_Vsel_0_(net1995[3]), .switch_n3_Vsel_1_(net1996[3]), .switch_n4_Vsel_0_(net1995[4]), .switch_n4_Vsel_1_(net1996[4]), .switch_n5_Vsel_0_(net1995[5]), .switch_n5_Vsel_1_(net1996[5]), .switch_n6_Vsel_0_(net1995[6]), .switch_n6_Vsel_1_(net1996[6]), .switch_n7_Vsel_0_(net2054[0]), .switch_n7_Vsel_1_(net2053[0]), .switch_n8_Vsel_0_(net2061[0]), .switch_n8_Vsel_1_(net2060[0]), .switch_n9_Vsel_0_(net2068[0]), .switch_n9_Vsel_1_(net2067[0]), .switch_n10_Vsel_0_(net2074[0]), .switch_n10_Vsel_1_(net2076[0]), .switch_n11_Vsel_0_(net2074[1]), .switch_n11_Vsel_1_(net2076[1]), .switch_n12_Vsel_0_(net2074[2]), .switch_n12_Vsel_1_(net2076[2]), .switch_n13_Vsel_0_(net2074[3]), .switch_n13_Vsel_1_(net2076[3]), .switch_n14_Vsel_0_(net2074[4]), .switch_n14_Vsel_1_(net2076[4]), .switch_n15_Vsel_0_(net2074[5]), .switch_n15_Vsel_1_(net2076[5]), .switch_n16_Vsel_0_(net2074[6]), .switch_n16_Vsel_1_(net2076[6]), .switch_n17_Vsel_0_(net2074[7]), .switch_n17_Vsel_1_(net2076[7]), .switch_n0_Vg_global_0_(net2009[0]), .switch_n0_Vg_global_1_(net2010[0]), .switch_n1_Vg_global_0_(net2009[1]), .switch_n1_Vg_global_1_(net2010[1]), .switch_n2_Vg_global_0_(net2009[2]), .switch_n2_Vg_global_1_(net2010[2]), .switch_n3_Vg_global_0_(net2009[3]), .switch_n3_Vg_global_1_(net2010[3]), .switch_n4_Vg_global_0_(net2009[4]), .switch_n4_Vg_global_1_(net2010[4]), .switch_n5_Vg_global_0_(net2009[5]), .switch_n5_Vg_global_1_(net2010[5]), .switch_n6_Vg_global_0_(net2009[6]), .switch_n6_Vg_global_1_(net2010[6]), .switch_n7_Vg_global_0_(net2056[0]), .switch_n7_Vg_global_1_(net2055[0]), .switch_n8_Vg_global_0_(net2063[0]), .switch_n8_Vg_global_1_(net2062[0]), .switch_n9_Vg_global_0_(net2070[0]), .switch_n9_Vg_global_1_(net2069[0]), .switch_n10_Vg_global_0_(net304[0]), .switch_n10_Vg_global_1_(net305[0]), .switch_n11_Vg_global_0_(net304[1]), .switch_n11_Vg_global_1_(net305[1]), .switch_n12_Vg_global_0_(net304[2]), .switch_n12_Vg_global_1_(net305[2]), .switch_n13_Vg_global_0_(net304[3]), .switch_n13_Vg_global_1_(net305[3]), .switch_n14_Vg_global_0_(net304[4]), .switch_n14_Vg_global_1_(net305[4]), .switch_n15_Vg_global_0_(net304[5]), .switch_n15_Vg_global_1_(net305[5]), .switch_n16_Vg_global_0_(net304[6]), .switch_n16_Vg_global_1_(net305[6]), .switch_n17_Vg_global_0_(net304[7]), .switch_n17_Vg_global_1_(net305[7]), .switch_n0_VTUN(net2023[0]), .switch_n1_VTUN(net2023[1]), .switch_n2_VTUN(net2023[2]), .switch_n3_VTUN(net2023[3]), .switch_n4_VTUN(net2023[4]), .switch_n5_VTUN(net2023[5]), .switch_n6_VTUN(net2023[6]), .switch_n7_VTUN(net2051[0]), .switch_n8_VTUN(net2058[0]), .switch_n9_VTUN(net2065[0]), .switch_n10_VTUN(net2071[0]), .switch_n11_VTUN(net2071[1]), .switch_n12_VTUN(net2071[2]), .switch_n13_VTUN(net2071[3]), .switch_n14_VTUN(net2071[4]), .switch_n15_VTUN(net2071[5]), .switch_n16_VTUN(net2071[6]), .switch_n17_VTUN(net2071[7]), .switch_n0_VINJ(net2037[0]), .switch_n1_VINJ(net2037[1]), .switch_n2_VINJ(net2037[2]), .switch_n3_VINJ(net2037[3]), .switch_n4_VINJ(net2037[4]), .switch_n5_VINJ(net2037[5]), .switch_n6_VINJ(net2037[6]), .switch_n7_VINJ(net2050[0]), .switch_n8_VINJ(net2057[0]), .switch_n9_VINJ(net2064[0]), .switch_n10_VINJ(net2072[0]), .switch_n11_VINJ(net2072[1]), .switch_n12_VINJ(net2072[2]), .switch_n13_VINJ(net2072[3]), .switch_n14_VINJ(net2072[4]), .switch_n15_VINJ(net2072[5]), .switch_n16_VINJ(net2072[6]), .switch_n17_VINJ(net2072[7]));
	none switch_ind(.island_num(1), .direction(horizontal), .col(18));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(19), .VPWR_0_(net1994), .VPWR_1_(net1994), .GND_T(net2073[8]), .VTUN_T(net2071[8]), .decode_0_(net2074[8]), .decode_1_(net2076[8]), .VINJ_T(net2072[8]), .GND(net1907), .CTRL_B_0_(net1972), .CTRL_B_1_(net1973), .run_r(net1903), .prog_r(net1904), .Vg_0_(net1974), .Vg_1_(net1975), .VTUN(net1905), .VINJ(net1906), .VDD_1_(net2317[0]));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net1148[0:6]), .out_1_row_0(net1149[0:6]), .VINJ_0_row_0(net1152[0:6]), .VINJ_1_row_0(net1153[0:6]), .Vsel_0_row_0(net1156[0:6]), .Vsel_1_row_0(net1157[0:6]), .Vg_0_row_0(net1160[0:6]), .Vg_1_row_0(net1161[0:6]), .GNDrow_0(net1138[0:6]), .VTUNrow_0(net1164[0:6]), .Dcol_0(net124[6:7]), .CLKcol_0(net125[6:7]), .Qcol_5(net125[6:7]), .comcol_0(net2316[0:1]), .VDDcol_0(net2317[0:1]), .Vd_Pcol_0(net2318[0:1]));
=======
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(1), .direction(vertical), .num(12), .type(prog_switch), .switch_n8_PR_0_(net2504[0]), .switch_n8_PR_1_(net2508[0]), .switch_n8_PR_2_(net2512[0]), .switch_n8_PR_3_(net2516[0]), .switch_n8_In_0_(net2503[0]), .switch_n8_In_1_(net2507[0]), .switch_n8_In_2_(net2511[0]), .switch_n8_In_3_(net2515[0]));
	TSMC350nm_GorS_IndrctSwcs switch(.island_num(1), .direction(horizontal), .num(20), .switch_n0_Input_0_(net2183), .switch_n0_Input_1_(net2219[0]), .switch_n1_Input_0_(net124[1]), .switch_n1_Input_1_(net125[1]), .switch_n2_Input_0_(net124[2]), .switch_n2_Input_1_(net125[2]), .switch_n3_Input_0_(net124[3]), .switch_n3_Input_1_(net125[3]), .switch_n4_Input_0_(net326[0]), .switch_n4_Input_1_(net327[0]), .switch_n5_Input_0_(net326[1]), .switch_n5_Input_1_(net327[1]), .switch_n6_Input_0_(net326[2]), .switch_n6_Input_1_(net327[2]), .switch_n7_Input_0_(net326[3]), .switch_n7_Input_1_(net327[3]), .switch_n8_Input_0_(net2502[0]), .switch_n8_Input_1_(net2089[0]), .switch_n9_Input_0_(net2090[0]), .switch_n9_Input_1_(net2102[0]), .switch_n10_Input_0_(net2103[0]), .switch_n10_Input_1_(net2120[0]), .switch_n11_Input_0_(net2121[0]), .switch_n11_Input_1_(net2140[0]), .switch_n12_Input_0_(net2141[0]), .switch_n12_Input_1_(net2142[0]), .switch_n13_Input_0_(net2143[0]), .switch_n13_Input_1_(net2144[0]), .switch_n14_Input_0_(net2145[0]), .switch_n14_Input_1_(net2157[0]), .switch_n15_Input_0_(net2158[0]), .switch_n15_Input_1_(net2170[0]), .switch_n16_Input_0_(net2171[0]), .switch_n16_Input_1_(net2178[0]), .switch_n17_Input_0_(net2179[0]), .switch_n17_Input_1_(net2180[0]), .switch_n0_GND(net2219[0]), .switch_n1_GND(net2219[1]), .switch_n2_GND(net2219[2]), .switch_n3_GND(net2219[3]), .switch_n4_GND(net2219[4]), .switch_n5_GND(net2219[5]), .switch_n6_GND(net2219[6]), .switch_n7_GND(net2241[0]), .switch_n8_GND(net2248[0]), .switch_n9_GND(net2255[0]), .switch_n10_GND(net325[0]), .switch_n11_GND(net325[1]), .switch_n12_GND(net325[2]), .switch_n13_GND(net325[3]), .switch_n14_GND(net325[4]), .switch_n15_GND(net325[5]), .switch_n16_GND(net325[6]), .switch_n17_GND(net325[7]), .switch_n0_Vsel_0_(net2184[0]), .switch_n0_Vsel_1_(net2185[0]), .switch_n1_Vsel_0_(net2184[1]), .switch_n1_Vsel_1_(net2185[1]), .switch_n2_Vsel_0_(net2184[2]), .switch_n2_Vsel_1_(net2185[2]), .switch_n3_Vsel_0_(net2184[3]), .switch_n3_Vsel_1_(net2185[3]), .switch_n4_Vsel_0_(net2184[4]), .switch_n4_Vsel_1_(net2185[4]), .switch_n5_Vsel_0_(net2184[5]), .switch_n5_Vsel_1_(net2185[5]), .switch_n6_Vsel_0_(net2184[6]), .switch_n6_Vsel_1_(net2185[6]), .switch_n7_Vsel_0_(net2243[0]), .switch_n7_Vsel_1_(net2242[0]), .switch_n8_Vsel_0_(net2250[0]), .switch_n8_Vsel_1_(net2249[0]), .switch_n9_Vsel_0_(net2257[0]), .switch_n9_Vsel_1_(net2256[0]), .switch_n10_Vsel_0_(net2263[0]), .switch_n10_Vsel_1_(net2265[0]), .switch_n11_Vsel_0_(net2263[1]), .switch_n11_Vsel_1_(net2265[1]), .switch_n12_Vsel_0_(net2263[2]), .switch_n12_Vsel_1_(net2265[2]), .switch_n13_Vsel_0_(net2263[3]), .switch_n13_Vsel_1_(net2265[3]), .switch_n14_Vsel_0_(net2263[4]), .switch_n14_Vsel_1_(net2265[4]), .switch_n15_Vsel_0_(net2263[5]), .switch_n15_Vsel_1_(net2265[5]), .switch_n16_Vsel_0_(net2263[6]), .switch_n16_Vsel_1_(net2265[6]), .switch_n17_Vsel_0_(net2263[7]), .switch_n17_Vsel_1_(net2265[7]), .switch_n0_Vg_global_0_(net2198[0]), .switch_n0_Vg_global_1_(net2199[0]), .switch_n1_Vg_global_0_(net2198[1]), .switch_n1_Vg_global_1_(net2199[1]), .switch_n2_Vg_global_0_(net2198[2]), .switch_n2_Vg_global_1_(net2199[2]), .switch_n3_Vg_global_0_(net2198[3]), .switch_n3_Vg_global_1_(net2199[3]), .switch_n4_Vg_global_0_(net2198[4]), .switch_n4_Vg_global_1_(net2199[4]), .switch_n5_Vg_global_0_(net2198[5]), .switch_n5_Vg_global_1_(net2199[5]), .switch_n6_Vg_global_0_(net2198[6]), .switch_n6_Vg_global_1_(net2199[6]), .switch_n7_Vg_global_0_(net2245[0]), .switch_n7_Vg_global_1_(net2244[0]), .switch_n8_Vg_global_0_(net2252[0]), .switch_n8_Vg_global_1_(net2251[0]), .switch_n9_Vg_global_0_(net2259[0]), .switch_n9_Vg_global_1_(net2258[0]), .switch_n10_Vg_global_0_(net346[0]), .switch_n10_Vg_global_1_(net347[0]), .switch_n11_Vg_global_0_(net346[1]), .switch_n11_Vg_global_1_(net347[1]), .switch_n12_Vg_global_0_(net346[2]), .switch_n12_Vg_global_1_(net347[2]), .switch_n13_Vg_global_0_(net346[3]), .switch_n13_Vg_global_1_(net347[3]), .switch_n14_Vg_global_0_(net346[4]), .switch_n14_Vg_global_1_(net347[4]), .switch_n15_Vg_global_0_(net346[5]), .switch_n15_Vg_global_1_(net347[5]), .switch_n16_Vg_global_0_(net346[6]), .switch_n16_Vg_global_1_(net347[6]), .switch_n17_Vg_global_0_(net346[7]), .switch_n17_Vg_global_1_(net347[7]), .switch_n0_VTUN(net2212[0]), .switch_n1_VTUN(net2212[1]), .switch_n2_VTUN(net2212[2]), .switch_n3_VTUN(net2212[3]), .switch_n4_VTUN(net2212[4]), .switch_n5_VTUN(net2212[5]), .switch_n6_VTUN(net2212[6]), .switch_n7_VTUN(net2240[0]), .switch_n8_VTUN(net2247[0]), .switch_n9_VTUN(net2254[0]), .switch_n10_VTUN(net348[0]), .switch_n11_VTUN(net348[1]), .switch_n12_VTUN(net348[2]), .switch_n13_VTUN(net348[3]), .switch_n14_VTUN(net348[4]), .switch_n15_VTUN(net348[5]), .switch_n16_VTUN(net348[6]), .switch_n17_VTUN(net348[7]), .switch_n0_VINJ(net2226[0]), .switch_n1_VINJ(net2226[1]), .switch_n2_VINJ(net2226[2]), .switch_n3_VINJ(net2226[3]), .switch_n4_VINJ(net2226[4]), .switch_n5_VINJ(net2226[5]), .switch_n6_VINJ(net2226[6]), .switch_n7_VINJ(net2239[0]), .switch_n8_VINJ(net2246[0]), .switch_n9_VINJ(net2253[0]), .switch_n10_VINJ(net345[0]), .switch_n11_VINJ(net345[1]), .switch_n12_VINJ(net345[2]), .switch_n13_VINJ(net345[3]), .switch_n14_VINJ(net345[4]), .switch_n15_VINJ(net345[5]), .switch_n16_VINJ(net345[6]), .switch_n17_VINJ(net345[7]));
	none switch_ind(.island_num(1), .direction(horizontal), .col(18));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(1), .direction(horizontal), .col(19), .VPWR_0_(net2183), .VPWR_1_(net2183), .decode_0_(net2263[8]), .decode_1_(net2265[8]), .GND(net2095), .CTRL_B_0_(net2160), .CTRL_B_1_(net2161), .run_r(net2091), .prog_r(net2092), .Vg_0_(net2162), .Vg_1_(net2163), .VTUN(net2093), .VINJ(net2094), .VDD_1_(net2172));


	/* Island 2 */
	TSMC350nm_volatile_swcs I__0 (.island_num(2), .row(0), .col(0), .matrix_row(1), .matrix_col(6), .out_0_row_0(net1231[0:6]), .out_1_row_0(net1232[0:6]), .VINJ_0_row_0(net1235[0:6]), .VINJ_1_row_0(net1236[0:6]), .Vsel_0_row_0(net1239[0:6]), .Vsel_1_row_0(net1240[0:6]), .Vg_0_row_0(net1243[0:6]), .Vg_1_row_0(net1244[0:6]), .GNDrow_0(net1221[0:6]), .VTUNrow_0(net1247[0:6]), .Dcol_0(net124[6:7]), .CLKcol_0(net125[6:7]), .Qcol_5(net125[6:7]), .comcol_0(net2502[0:1]), .Vd_Pcol_0(net2516[0:1]), .Vd_in_0_col_0(net2503[0:1]), .Vd_in_1_col_0(net2507[0:1]), .Vd_in_2_col_0(net2511[0:1]), .Vd_in_3_col_0(net2515[0:1]), .Vd_in_4_col_0(net2504[0:1]), .Vd_in_5_col_0(net2508[0:1]), .Vd_in_6_col_0(net2512[0:1]), .Vd_in_7_col_0(net2516[0:1]), .Vd_o_0_col_5(net1917[0:1]), .Vd_o_1_col_5(net1918[0:1]), .Vd_o_2_col_5(net1919[0:1]), .Vd_o_3_col_5(net1920[0:1]), .Vd_o_4_col_5(net1921[0:1]), .Vd_o_5_col_5(net1922[0:1]), .Vd_o_6_col_5(net1923[0:1]), .Vd_o_7_col_5(net1924[0:1]));
>>>>>>> Stashed changes

 	/*Programming Mux */ 

 endmodule